module sram (
	// inout  wire [15:0]	dq
    // output wire [17:0]	addr
    // output wire 		ub_n
    // output wire 		lb_n
    // output wire 		we_n
    // output wire 		ce_n
    // output wire 		oe_n
);

endmodule
