// megafunction wizard: %Serial Flash Loader%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: altserial_flash_loader 

// ============================================================
// File Name: sfl.v
// Megafunction Name(s):
// 			altserial_flash_loader
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sfl (
	noe_in);

	input	  noe_in;


	altserial_flash_loader	altserial_flash_loader_component (
				.noe (noe_in)
				// synopsys translate_off
				,
				.asmi_access_granted (),
				.asmi_access_request (),
				.data0out (),
				.data_in (),
				.data_oe (),
				.data_out (),
				.dclkin (),
				.scein (),
				.sdoin ()
				// synopsys translate_on
				);
	defparam
		altserial_flash_loader_component.enable_quad_spi_support = 0,
		altserial_flash_loader_component.enable_shared_access = "OFF",
		altserial_flash_loader_component.enhanced_mode = 1,
		altserial_flash_loader_component.intended_device_family = "Cyclone II";


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: ENABLE_QUAD_SPI_SUPPORT NUMERIC "0"
// Retrieval info: CONSTANT: ENABLE_SHARED_ACCESS STRING "OFF"
// Retrieval info: CONSTANT: ENHANCED_MODE NUMERIC "1"
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: USED_PORT: noe_in 0 0 0 0 INPUT NODEFVAL "noe_in"
// Retrieval info: CONNECT: @noe 0 0 0 0 noe_in 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL sfl.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sfl.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sfl.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sfl.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sfl_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sfl_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
