---------------------------------------------------------------------
-- File Name: filtebank_package.vhd
-- Module: filterbank
-- Function Description:
--	This module contains the constants and types and function
--	used by filterbank.vhd module. 
---------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_SIGNED.all;
use work.mul.all;

package filterbank_package is

constant MAX_OUTPUT_LIMIT	: integer := 32767;


type samples_type is array(0 to 31) of std_logic_vector(31 downto 0);
type pre_gen_return_type is array(0 to 31) of integer;

type table_D_type is array(0 to 511) of integer;
constant D : table_D_type := (
0 ,      -- 0.0000000000 */ ,
-16384 ,      -- -0.0000152590 */ ,
-16384 ,      -- -0.0000152590 */ ,
-16384 ,      -- -0.0000152590 */ ,
-16384 ,      -- -0.0000152590 */ ,
-16384 ,      -- -0.0000152590 */ ,
-16384 ,      -- -0.0000152590 */ ,
-32768 ,      -- -0.0000305180 */ ,
-32768 ,      -- -0.0000305180 */ ,
-32768 ,      -- -0.0000305180 */ ,
-32768 ,      -- -0.0000305180 */ ,
-49151 ,      -- -0.0000457760 */ ,
-49151 ,      -- -0.0000457760 */ ,
-65535 ,      -- -0.0000610350 */ ,
-65535 ,      -- -0.0000610350 */ ,
-81920 ,      -- -0.0000762940 */ ,
-81920 ,      -- -0.0000762940 */ ,
-98304 ,      -- -0.0000915530 */ ,
-114688 ,      -- -0.0001068120 */ ,
-114688 ,      -- -0.0001068120 */ ,
-131071 ,      -- -0.0001220700 */ ,
-147455 ,      -- -0.0001373290 */ ,
-163840 ,      -- -0.0001525880 */ ,
-180224 ,      -- -0.0001678470 */ ,
-212991 ,      -- -0.0001983640 */ ,
-229375 ,      -- -0.0002136230 */ ,
-262144 ,      -- -0.0002441410 */ ,
-278527 ,      -- -0.0002593990 */ ,
-311296 ,      -- -0.0002899170 */ ,
-344064 ,      -- -0.0003204350 */ ,
-393216 ,      -- -0.0003662110 */ ,
-425984 ,      -- -0.0003967290 */ ,
-475136 ,      -- -0.0004425050 */ ,
-507903 ,      -- -0.0004730220 */ ,
-573440 ,      -- -0.0005340580 */ ,
-622592 ,      -- -0.0005798340 */ ,
-671743 ,      -- -0.0006256100 */ ,
-737280 ,      -- -0.0006866460 */ ,
-802816 ,      -- -0.0007476810 */ ,
-868352 ,      -- -0.0008087160 */ ,
-950272 ,      -- -0.0008850100 */ ,
-1032192 ,      -- -0.0009613040 */ ,
-1114112 ,      -- -0.0010375980 */ ,
-1196032 ,      -- -0.0011138920 */ ,
-1294335 ,      -- -0.0012054440 */ ,
-1392639 ,      -- -0.0012969970 */ ,
-1490944 ,      -- -0.0013885500 */ ,
-1589248 ,      -- -0.0014801030 */ ,
-1703935 ,      -- -0.0015869140 */ ,
-1818624 ,      -- -0.0016937260 */ ,
-1916927 ,      -- -0.0017852780 */ ,
-2048000 ,      -- -0.0019073490 */ ,
-2162687 ,      -- -0.0020141600 */ ,
-2277376 ,      -- -0.0021209720 */ ,
-2408448 ,      -- -0.0022430420 */ ,
-2523136 ,      -- -0.0023498540 */ ,
-2637823 ,      -- -0.0024566650 */ ,
-2768895 ,      -- -0.0025787350 */ ,
-2883584 ,      -- -0.0026855470 */ ,
-2998271 ,      -- -0.0027923580 */ ,
-3112960 ,      -- -0.0028991700 */ ,
-3211264 ,      -- -0.0029907230 */ ,
-3309567 ,      -- -0.0030822750 */ ,
-3407871 ,      -- -0.0031738280 */ ,
3489791 ,      -- 0.0032501220 */ ,
3571711 ,      -- 0.0033264160 */ ,
3637247 ,      -- 0.0033874510 */ ,
3686400 ,      -- 0.0034332280 */ ,
3719167 ,      -- 0.0034637450 */ ,
3735552 ,      -- 0.0034790040 */ ,
3735552 ,      -- 0.0034790040 */ ,
3719167 ,      -- 0.0034637450 */ ,
3670016 ,      -- 0.0034179690 */ ,
3620863 ,      -- 0.0033721920 */ ,
3522560 ,      -- 0.0032806400 */ ,
3407871 ,      -- 0.0031738280 */ ,
3276800 ,      -- 0.0030517580 */ ,
3096575 ,      -- 0.0028839110 */ ,
2899968 ,      -- 0.0027008060 */ ,
2670592 ,      -- 0.0024871830 */ ,
2392063 ,      -- 0.0022277830 */ ,
2080767 ,      -- 0.0019378660 */ ,
1736704 ,      -- 0.0016174320 */ ,
1359871 ,      -- 0.0012664790 */ ,
933888 ,      -- 0.0008697510 */ ,
475136 ,      -- 0.0004425050 */ ,
-32768 ,      -- -0.0000305180 */ ,
-589823 ,      -- -0.0005493160 */ ,
-1179648 ,      -- -0.0010986330 */ ,
-1818624 ,      -- -0.0016937260 */ ,
-2506752 ,      -- -0.0023345950 */ ,
-3227647 ,      -- -0.0030059810 */ ,
-3997696 ,      -- -0.0037231450 */ ,
-4816896 ,      -- -0.0044860840 */ ,
-5685248 ,      -- -0.0052948000 */ ,
-6569983 ,      -- -0.0061187740 */ ,
-7520255 ,      -- -0.0070037840 */ ,
-8503296 ,      -- -0.0079193120 */ ,
-9519103 ,      -- -0.0088653560 */ ,
-10567680 ,      -- -0.0098419190 */ ,
-11649023 ,      -- -0.0108489990 */ ,
-12763136 ,      -- -0.0118865970 */ ,
-13893631 ,      -- -0.0129394530 */ ,
-15056895 ,      -- -0.0140228270 */ ,
-16236544 ,      -- -0.0151214600 */ ,
-17432576 ,      -- -0.0162353520 */ ,
-18628607 ,      -- -0.0173492430 */ ,
-19824640 ,      -- -0.0184631350 */ ,
-21020671 ,      -- -0.0195770260 */ ,
-22216704 ,      -- -0.0206909180 */ ,
-23396352 ,      -- -0.0217895510 */ ,
-24543231 ,      -- -0.0228576660 */ ,
-25673727 ,      -- -0.0239105220 */ ,
-26771455 ,      -- -0.0249328610 */ ,
-27820032 ,      -- -0.0259094240 */ ,
-28819456 ,      -- -0.0268402100 */ ,
-29769728 ,      -- -0.0277252200 */ ,
-30638080 ,      -- -0.0285339360 */ ,
-31440895 ,      -- -0.0292816160 */ ,
-32145407 ,      -- -0.0299377440 */ ,
-32784384 ,      -- -0.0305328370 */ ,
-33292287 ,      -- -0.0310058590 */ ,
-33701887 ,      -- -0.0313873290 */ ,
-33996799 ,      -- -0.0316619870 */ ,
-34160639 ,      -- -0.0318145750 */ ,
-34193408 ,      -- -0.0318450930 */ ,
-34078719 ,      -- -0.0317382810 */ ,
-33800192 ,      -- -0.0314788820 */ ,
33374207 ,      -- 0.0310821530 */ ,
32767999 ,      -- 0.0305175780 */ ,
31981567 ,      -- 0.0297851560 */ ,
31014912 ,      -- 0.0288848880 */ ,
29851648 ,      -- 0.0278015140 */ ,
28491775 ,      -- 0.0265350340 */ ,
26935295 ,      -- 0.0250854490 */ ,
25149439 ,      -- 0.0234222410 */ ,
23166976 ,      -- 0.0215759280 */ ,
20971520 ,      -- 0.0195312500 */ ,
18530303 ,      -- 0.0172576900 */ ,
15892479 ,      -- 0.0148010250 */ ,
13008896 ,      -- 0.0121154790 */ ,
9912319 ,      -- 0.0092315670 */ ,
6586367 ,      -- 0.0061340330 */ ,
3031040 ,      -- 0.0028228760 */ ,
-737280 ,      -- -0.0006866460 */ ,
-4718591 ,      -- -0.0043945310 */ ,
-8929279 ,      -- -0.0083160400 */ ,
-13336575 ,      -- -0.0124206540 */ ,
-17940479 ,      -- -0.0167083740 */ ,
-22740991 ,      -- -0.0211791990 */ ,
-27721727 ,      -- -0.0258178710 */ ,
-32866304 ,      -- -0.0306091310 */ ,
-38174720 ,      -- -0.0355529790 */ ,
-43630591 ,      -- -0.0406341550 */ ,
-49217535 ,      -- -0.0458374020 */ ,
-54902783 ,      -- -0.0511322020 */ ,
-60702719 ,      -- -0.0565338130 */ ,
-66568192 ,      -- -0.0619964600 */ ,
-72499200 ,      -- -0.0675201420 */ ,
-78446591 ,      -- -0.0730590820 */ ,
-84426751 ,      -- -0.0786285400 */ ,
-90390527 ,      -- -0.0841827390 */ ,
-96321536 ,      -- -0.0897064210 */ ,
-102187007 ,      -- -0.0951690670 */ ,
-107954175 ,      -- -0.1005401610 */ ,
-113623039 ,      -- -0.1058197020 */ ,
-119128063 ,      -- -0.1109466550 */ ,
-124469248 ,      -- -0.1159210210 */ ,
-129597439 ,      -- -0.1206970210 */ ,
-134496255 ,      -- -0.1252593990 */ ,
-139116544 ,      -- -0.1295623780 */ ,
-143441919 ,      -- -0.1335906980 */ ,
-147423232 ,      -- -0.1372985840 */ ,
-151044095 ,      -- -0.1406707760 */ ,
-154271744 ,      -- -0.1436767580 */ ,
-157040639 ,      -- -0.1462554930 */ ,
-159367167 ,      -- -0.1484222410 */ ,
-161185792 ,      -- -0.1501159670 */ ,
-162463743 ,      -- -0.1513061520 */ ,
-163168255 ,      -- -0.1519622800 */ ,
-163282944 ,      -- -0.1520690920 */ ,
-162775039 ,      -- -0.1515960690 */ ,
-161595392 ,      -- -0.1504974370 */ ,
-159743999 ,      -- -0.1487731930 */ ,
-157155328 ,      -- -0.1463623050 */ ,
-153829376 ,      -- -0.1432647710 */ ,
-149733375 ,      -- -0.1394500730 */ ,
-144834559 ,      -- -0.1348876950 */ ,
-139132928 ,      -- -0.1295776370 */ ,
-132579327 ,      -- -0.1234741210 */ ,
-125173759 ,      -- -0.1165771480 */ ,
-116883455 ,      -- -0.1088562010 */ ,
107708415 ,      -- 0.1003112790 */ ,
97632255 ,      -- 0.0909271240 */ ,
86638592 ,      -- 0.0806884770 */ ,
74727424 ,      -- 0.0695953370 */ ,
61865983 ,      -- 0.0576171870 */ ,
48087040 ,      -- 0.0447845460 */ ,
33374207 ,      -- 0.0310821530 */ ,
17727488 ,      -- 0.0165100100 */ ,
1146879 ,      -- 0.0010681150 */ ,
-16351231 ,      -- -0.0152282710 */ ,
-34766847 ,      -- -0.0323791500 */ ,
-54067200 ,      -- -0.0503540040 */ ,
-74268672 ,      -- -0.0691680910 */ ,
-95322112 ,      -- -0.0887756350 */ ,
-117211136 ,      -- -0.1091613770 */ ,
-139919360 ,      -- -0.1303100590 */ ,
-163430400 ,      -- -0.1522064210 */ ,
-187678720 ,      -- -0.1747894290 */ ,
-212664319 ,      -- -0.1980590820 */ ,
-238354431 ,      -- -0.2219848630 */ ,
-264683519 ,      -- -0.2465057370 */ ,
-291618816 ,      -- -0.2715911870 */ ,
-319127551 ,      -- -0.2972106930 */ ,
-347160575 ,      -- -0.3233184810 */ ,
-375668735 ,      -- -0.3498687740 */ ,
-404586495 ,      -- -0.3768005370 */ ,
-433881088 ,      -- -0.4040832520 */ ,
-463486976 ,      -- -0.4316558840 */ ,
-493355007 ,      -- -0.4594726560 */ ,
-523419647 ,      -- -0.4874725340 */ ,
-553631743 ,      -- -0.5156097410 */ ,
-583925759 ,      -- -0.5438232420 */ ,
-614219775 ,      -- -0.5720367430 */ ,
-644481024 ,      -- -0.6002197270 */ ,
-674627583 ,      -- -0.6282958980 */ ,
-704610303 ,      -- -0.6562194820 */ ,
-734347264 ,      -- -0.6839141850 */ ,
-763772928 ,      -- -0.7113189700 */ ,
-792821760 ,      -- -0.7383728030 */ ,
-821444607 ,      -- -0.7650299070 */ ,
-849559551 ,      -- -0.7912139890 */ ,
-877101056 ,      -- -0.8168640140 */ ,
-904036352 ,      -- -0.8419494630 */ ,
-930250751 ,      -- -0.8663635250 */ ,
-955727871 ,      -- -0.8900909420 */ ,
-980385792 ,      -- -0.9130554200 */ ,
-1004158976 ,      -- -0.9351959230 */ ,
-1027014656 ,      -- -0.9564819340 */ ,
-1048887296 ,      -- -0.9768524170 */ ,
-1069711360 ,      -- -0.9962463380 */ ,
-1089437696 ,      -- -1.0146179200 */ ,
-1108033536 ,      -- -1.0319366460 */ ,
-1125449727 ,      -- -1.0481567380 */ ,
-1141620735 ,      -- -1.0632171630 */ ,
-1156546560 ,      -- -1.0771179200 */ ,
-1170145280 ,      -- -1.0897827150 */ ,
-1182416896 ,      -- -1.1012115480 */ ,
-1193328639 ,      -- -1.1113739010 */ ,
-1202831359 ,      -- -1.1202239990 */ ,
-1210908671 ,      -- -1.1277465820 */ ,
-1217544192 ,      -- -1.1339263920 */ ,
-1222737920 ,      -- -1.1387634280 */ ,
-1226440703 ,      -- -1.1422119140 */ ,
-1228668927 ,      -- -1.1442871090 */ ,
1229422592 ,      -- 1.1449890140 */ ,
1228668927 ,      -- 1.1442871090 */ ,
1226440703 ,      -- 1.1422119140 */ ,
1222737920 ,      -- 1.1387634280 */ ,
1217544192 ,      -- 1.1339263920 */ ,
1210908671 ,      -- 1.1277465820 */ ,
1202831359 ,      -- 1.1202239990 */ ,
1193328639 ,      -- 1.1113739010 */ ,
1182416896 ,      -- 1.1012115480 */ ,
1170145280 ,      -- 1.0897827150 */ ,
1156546560 ,      -- 1.0771179200 */ ,
1141620735 ,      -- 1.0632171630 */ ,
1125449727 ,      -- 1.0481567380 */ ,
1108033536 ,      -- 1.0319366460 */ ,
1089437696 ,      -- 1.0146179200 */ ,
1069711360 ,      -- 0.9962463380 */ ,
1048887296 ,      -- 0.9768524170 */ ,
1027014656 ,      -- 0.9564819340 */ ,
1004158976 ,      -- 0.9351959230 */ ,
980385792 ,      -- 0.9130554200 */ ,
955727871 ,      -- 0.8900909420 */ ,
930250751 ,      -- 0.8663635250 */ ,
904036352 ,      -- 0.8419494630 */ ,
877101056 ,      -- 0.8168640140 */ ,
849559551 ,      -- 0.7912139890 */ ,
821444607 ,      -- 0.7650299070 */ ,
792821760 ,      -- 0.7383728030 */ ,
763772928 ,      -- 0.7113189700 */ ,
734347264 ,      -- 0.6839141850 */ ,
704610303 ,      -- 0.6562194820 */ ,
674627583 ,      -- 0.6282958980 */ ,
644481024 ,      -- 0.6002197270 */ ,
614219775 ,      -- 0.5720367430 */ ,
583925759 ,      -- 0.5438232420 */ ,
553631743 ,      -- 0.5156097410 */ ,
523419647 ,      -- 0.4874725340 */ ,
493355007 ,      -- 0.4594726560 */ ,
463486976 ,      -- 0.4316558840 */ ,
433881088 ,      -- 0.4040832520 */ ,
404586495 ,      -- 0.3768005370 */ ,
375668735 ,      -- 0.3498687740 */ ,
347160575 ,      -- 0.3233184810 */ ,
319127551 ,      -- 0.2972106930 */ ,
291618816 ,      -- 0.2715911870 */ ,
264683519 ,      -- 0.2465057370 */ ,
238354431 ,      -- 0.2219848630 */ ,
212664319 ,      -- 0.1980590820 */ ,
187678720 ,      -- 0.1747894290 */ ,
163430400 ,      -- 0.1522064210 */ ,
139919360 ,      -- 0.1303100590 */ ,
117211136 ,      -- 0.1091613770 */ ,
95322112 ,      -- 0.0887756350 */ ,
74268672 ,      -- 0.0691680910 */ ,
54067200 ,      -- 0.0503540040 */ ,
34766847 ,      -- 0.0323791500 */ ,
16351231 ,      -- 0.0152282710 */ ,
-1146879 ,      -- -0.0010681150 */ ,
-17727488 ,      -- -0.0165100100 */ ,
-33374207 ,      -- -0.0310821530 */ ,
-48087040 ,      -- -0.0447845460 */ ,
-61865983 ,      -- -0.0576171870 */ ,
-74727424 ,      -- -0.0695953370 */ ,
-86638592 ,      -- -0.0806884770 */ ,
-97632255 ,      -- -0.0909271240 */ ,
107708415 ,      -- 0.1003112790 */ ,
116883455 ,      -- 0.1088562010 */ ,
125173759 ,      -- 0.1165771480 */ ,
132579327 ,      -- 0.1234741210 */ ,
139132928 ,      -- 0.1295776370 */ ,
144834559 ,      -- 0.1348876950 */ ,
149733375 ,      -- 0.1394500730 */ ,
153829376 ,      -- 0.1432647710 */ ,
157155328 ,      -- 0.1463623050 */ ,
159743999 ,      -- 0.1487731930 */ ,
161595392 ,      -- 0.1504974370 */ ,
162775039 ,      -- 0.1515960690 */ ,
163282944 ,      -- 0.1520690920 */ ,
163168255 ,      -- 0.1519622800 */ ,
162463743 ,      -- 0.1513061520 */ ,
161185792 ,      -- 0.1501159670 */ ,
159367167 ,      -- 0.1484222410 */ ,
157040639 ,      -- 0.1462554930 */ ,
154271744 ,      -- 0.1436767580 */ ,
151044095 ,      -- 0.1406707760 */ ,
147423232 ,      -- 0.1372985840 */ ,
143441919 ,      -- 0.1335906980 */ ,
139116544 ,      -- 0.1295623780 */ ,
134496255 ,      -- 0.1252593990 */ ,
129597439 ,      -- 0.1206970210 */ ,
124469248 ,      -- 0.1159210210 */ ,
119128063 ,      -- 0.1109466550 */ ,
113623039 ,      -- 0.1058197020 */ ,
107954175 ,      -- 0.1005401610 */ ,
102187007 ,      -- 0.0951690670 */ ,
96321536 ,      -- 0.0897064210 */ ,
90390527 ,      -- 0.0841827390 */ ,
84426751 ,      -- 0.0786285400 */ ,
78446591 ,      -- 0.0730590820 */ ,
72499200 ,      -- 0.0675201420 */ ,
66568192 ,      -- 0.0619964600 */ ,
60702719 ,      -- 0.0565338130 */ ,
54902783 ,      -- 0.0511322020 */ ,
49217535 ,      -- 0.0458374020 */ ,
43630591 ,      -- 0.0406341550 */ ,
38174720 ,      -- 0.0355529790 */ ,
32866304 ,      -- 0.0306091310 */ ,
27721727 ,      -- 0.0258178710 */ ,
22740991 ,      -- 0.0211791990 */ ,
17940479 ,      -- 0.0167083740 */ ,
13336575 ,      -- 0.0124206540 */ ,
8929279 ,      -- 0.0083160400 */ ,
4718591 ,      -- 0.0043945310 */ ,
737280 ,      -- 0.0006866460 */ ,
-3031040 ,      -- -0.0028228760 */ ,
-6586367 ,      -- -0.0061340330 */ ,
-9912319 ,      -- -0.0092315670 */ ,
-13008896 ,      -- -0.0121154790 */ ,
-15892479 ,      -- -0.0148010250 */ ,
-18530303 ,      -- -0.0172576900 */ ,
-20971520 ,      -- -0.0195312500 */ ,
-23166976 ,      -- -0.0215759280 */ ,
-25149439 ,      -- -0.0234222410 */ ,
-26935295 ,      -- -0.0250854490 */ ,
-28491775 ,      -- -0.0265350340 */ ,
-29851648 ,      -- -0.0278015140 */ ,
-31014912 ,      -- -0.0288848880 */ ,
-31981567 ,      -- -0.0297851560 */ ,
-32767999 ,      -- -0.0305175780 */ ,
33374207 ,      -- 0.0310821530 */ ,
33800192 ,      -- 0.0314788820 */ ,
34078719 ,      -- 0.0317382810 */ ,
34193408 ,      -- 0.0318450930 */ ,
34160639 ,      -- 0.0318145750 */ ,
33996799 ,      -- 0.0316619870 */ ,
33701887 ,      -- 0.0313873290 */ ,
33292287 ,      -- 0.0310058590 */ ,
32784384 ,      -- 0.0305328370 */ ,
32145407 ,      -- 0.0299377440 */ ,
31440895 ,      -- 0.0292816160 */ ,
30638080 ,      -- 0.0285339360 */ ,
29769728 ,      -- 0.0277252200 */ ,
28819456 ,      -- 0.0268402100 */ ,
27820032 ,      -- 0.0259094240 */ ,
26771455 ,      -- 0.0249328610 */ ,
25673727 ,      -- 0.0239105220 */ ,
24543231 ,      -- 0.0228576660 */ ,
23396352 ,      -- 0.0217895510 */ ,
22216704 ,      -- 0.0206909180 */ ,
21020671 ,      -- 0.0195770260 */ ,
19824640 ,      -- 0.0184631350 */ ,
18628607 ,      -- 0.0173492430 */ ,
17432576 ,      -- 0.0162353520 */ ,
16236544 ,      -- 0.0151214600 */ ,
15056895 ,      -- 0.0140228270 */ ,
13893631 ,      -- 0.0129394530 */ ,
12763136 ,      -- 0.0118865970 */ ,
11649023 ,      -- 0.0108489990 */ ,
10567680 ,      -- 0.0098419190 */ ,
9519103 ,      -- 0.0088653560 */ ,
8503296 ,      -- 0.0079193120 */ ,
7520255 ,      -- 0.0070037840 */ ,
6569983 ,      -- 0.0061187740 */ ,
5685248 ,      -- 0.0052948000 */ ,
4816896 ,      -- 0.0044860840 */ ,
3997696 ,      -- 0.0037231450 */ ,
3227647 ,      -- 0.0030059810 */ ,
2506752 ,      -- 0.0023345950 */ ,
1818624 ,      -- 0.0016937260 */ ,
1179648 ,      -- 0.0010986330 */ ,
589823 ,      -- 0.0005493160 */ ,
32768 ,      -- 0.0000305180 */ ,
-475136 ,      -- -0.0004425050 */ ,
-933888 ,      -- -0.0008697510 */ ,
-1359871 ,      -- -0.0012664790 */ ,
-1736704 ,      -- -0.0016174320 */ ,
-2080767 ,      -- -0.0019378660 */ ,
-2392063 ,      -- -0.0022277830 */ ,
-2670592 ,      -- -0.0024871830 */ ,
-2899968 ,      -- -0.0027008060 */ ,
-3096575 ,      -- -0.0028839110 */ ,
-3276800 ,      -- -0.0030517580 */ ,
-3407871 ,      -- -0.0031738280 */ ,
-3522560 ,      -- -0.0032806400 */ ,
-3620863 ,      -- -0.0033721920 */ ,
-3670016 ,      -- -0.0034179690 */ ,
-3719167 ,      -- -0.0034637450 */ ,
-3735552 ,      -- -0.0034790040 */ ,
-3735552 ,      -- -0.0034790040 */ ,
-3719167 ,      -- -0.0034637450 */ ,
-3686400 ,      -- -0.0034332280 */ ,
-3637247 ,      -- -0.0033874510 */ ,
-3571711 ,      -- -0.0033264160 */ ,
3489791 ,      -- 0.0032501220 */ ,
3407871 ,      -- 0.0031738280 */ ,
3309567 ,      -- 0.0030822750 */ ,
3211264 ,      -- 0.0029907230 */ ,
3112960 ,      -- 0.0028991700 */ ,
2998271 ,      -- 0.0027923580 */ ,
2883584 ,      -- 0.0026855470 */ ,
2768895 ,      -- 0.0025787350 */ ,
2637823 ,      -- 0.0024566650 */ ,
2523136 ,      -- 0.0023498540 */ ,
2408448 ,      -- 0.0022430420 */ ,
2277376 ,      -- 0.0021209720 */ ,
2162687 ,      -- 0.0020141600 */ ,
2048000 ,      -- 0.0019073490 */ ,
1916927 ,      -- 0.0017852780 */ ,
1818624 ,      -- 0.0016937260 */ ,
1703935 ,      -- 0.0015869140 */ ,
1589248 ,      -- 0.0014801030 */ ,
1490944 ,      -- 0.0013885500 */ ,
1392639 ,      -- 0.0012969970 */ ,
1294335 ,      -- 0.0012054440 */ ,
1196032 ,      -- 0.0011138920 */ ,
1114112 ,      -- 0.0010375980 */ ,
1032192 ,      -- 0.0009613040 */ ,
950272 ,      -- 0.0008850100 */ ,
868352 ,      -- 0.0008087160 */ ,
802816 ,      -- 0.0007476810 */ ,
737280 ,      -- 0.0006866460 */ ,
671743 ,      -- 0.0006256100 */ ,
622592 ,      -- 0.0005798340 */ ,
573440 ,      -- 0.0005340580 */ ,
507903 ,      -- 0.0004730220 */ ,
475136 ,      -- 0.0004425050 */ ,
425984 ,      -- 0.0003967290 */ ,
393216 ,      -- 0.0003662110 */ ,
344064 ,      -- 0.0003204350 */ ,
311296 ,      -- 0.0002899170 */ ,
278527 ,      -- 0.0002593990 */ ,
262144 ,      -- 0.0002441410 */ ,
229375 ,      -- 0.0002136230 */ ,
212991 ,      -- 0.0001983640 */ ,
180224 ,      -- 0.0001678470 */ ,
163840 ,      -- 0.0001525880 */ ,
147455 ,      -- 0.0001373290 */ ,
131071 ,      -- 0.0001220700 */ ,
114688 ,      -- 0.0001068120 */ ,
114688 ,      -- 0.0001068120 */ ,
98304 ,      -- 0.0000915530 */ ,
81920 ,      -- 0.0000762940 */ ,
81920 ,      -- 0.0000762940 */ ,
65535 ,      -- 0.0000610350 */ ,
65535 ,      -- 0.0000610350 */ ,
49151 ,      -- 0.0000457760 */ ,
49151 ,      -- 0.0000457760 */ ,
32768 ,      -- 0.0000305180 */ ,
32768 ,      -- 0.0000305180 */ ,
32768 ,      -- 0.0000305180 */ ,
32768 ,      -- 0.0000305180 */ ,
16384 ,      -- 0.0000152590 */ ,
16384 ,      -- 0.0000152590 */ ,
16384 ,      -- 0.0000152590 */ ,
16384 ,      -- 0.0000152590 */ ,
16384 ,      -- 0.0000152590 */ ,
16384 );      -- 0.0000152590 */


function subsyn_pre_gen(bandPtr_fix: samples_type; v_offset : integer ) return pre_gen_return_type;



end;



package body filterbank_package is

   function subsyn_pre_gen(bandPtr_fix: samples_type; v_offset : integer ) return pre_gen_return_type is
      type t_type is array(0 to 49) of integer;
      variable t : t_type;
      
      variable VOffsetPtr : pre_gen_return_type ;
   begin
        t(0) := conv_integer(bandPtr_fix(21));
	t(1) := conv_integer(bandPtr_fix(20));
	t(2) := conv_integer(bandPtr_fix(22));
	t(3) := conv_integer(bandPtr_fix(23));
	t(4) := conv_integer(bandPtr_fix(18));
	t(5) := conv_integer(bandPtr_fix(19));
	t(6) := conv_integer(bandPtr_fix(17));
	t(7) := conv_integer(bandPtr_fix(16));
	t(8) := conv_integer(bandPtr_fix(26));
	t(9) := conv_integer(bandPtr_fix(27));
	t(10) := conv_integer(bandPtr_fix(25));
	t(11) := conv_integer(bandPtr_fix(24));
	t(12) := conv_integer(bandPtr_fix(29));
	t(13) := conv_integer(bandPtr_fix(28));
	t(14) := conv_integer(bandPtr_fix(30));
	t(15) := conv_integer(bandPtr_fix(31));
	t(16) := conv_integer(bandPtr_fix(10));
	t(17) := conv_integer(bandPtr_fix(11));
	t(18) := conv_integer(bandPtr_fix(9));
	t(19) := conv_integer(bandPtr_fix(8));
	t(20) := conv_integer(bandPtr_fix(13));
	t(21) := conv_integer(bandPtr_fix(12));
	t(22) := conv_integer(bandPtr_fix(14));
	t(23) := conv_integer(bandPtr_fix(15));
	t(24) := conv_integer(bandPtr_fix(5));
	t(25) := conv_integer(bandPtr_fix(4));
	t(26) := conv_integer(bandPtr_fix(6));
	t(27) := conv_integer(bandPtr_fix(7));
	t(28) := conv_integer(bandPtr_fix(2));
	t(29) := conv_integer(bandPtr_fix(3));
	t(30) := conv_integer(bandPtr_fix(1));
	t(31) := conv_integer(bandPtr_fix(0));
	t(32) := t(16) + t(0);
	t(33) := t(16) - t(0);
	t(0) := fix_mul(1044287193, t(33));
	t(16) := t(17) + t(1);
	t(33) := t(17) - t(1);
	t(1) := fix_mul(627838283, t(33)) * 2;
	t(17) := t(18) + t(2);
	t(33) := t(18) - t(2);
	t(2) := fix_mul(901244819, t(33));
	t(18) := t(19) + t(3);
	t(33) := t(19) - t(3);
	t(3) := fix_mul(799439733, t(33));
	t(19) := t(20) + t(4);
	t(33) := t(20) - t(4);
	t(4) := fix_mul(552381383, t(33)) * 4;
	t(20) := t(21) + t(5);
	t(33) := t(21) - t(5);
	t(5) := fix_mul(796804811, t(33)) * 2;
	t(21) := t(22) + t(6);
	t(33) := t(22) - t(6);
	t(6) := fix_mul(914722919, t(33)) * 4;
	t(22) := t(23) + t(7);
	t(33) := t(23) - t(7);
	t(7) := fix_mul(683839869, t(33)) * 16;
	t(23) := t(24) + t(8);
	t(33) := t(24) - t(8);
	t(8) := fix_mul(625921656, t(33));
	t(24) := t(25) + t(9);
	t(33) := t(25) - t(9);
	t(9) := fix_mul(593890786, t(33));
	t(25) := t(26) + t(10);
	t(33) := t(26) - t(10);
	t(10) := fix_mul(668408712, t(33));
	t(26) := t(27) + t(11);
	t(33) := t(27) - t(11);
	t(11) := fix_mul(724569939, t(33));
	t(27) := t(28) + t(12);
	t(33) := t(28) - t(12);
	t(12) := fix_mul(553457334, t(33));
	t(28) := t(29) + t(13);
	t(33) := t(29) - t(13);
	t(13) := fix_mul(570202640, t(33));
	t(29) := t(30) + t(14);
	t(33) := t(30) - t(14);
	t(14) := fix_mul(542745310, t(33));
	t(30) := t(31) + t(15);
	t(33) := t(31) - t(15);
	t(15) := fix_mul(537518376, t(33));
	t(31) := t(8) + t(0);
	t(33) := t(8) - t(0);
	t(0) := fix_mul(569446996, t(33)) * 2;
	t(8) := t(9) + t(1);
	t(33) := t(9) - t(1);
	t(1) := fix_mul(846274582, t(33));
	t(9) := t(10) + t(2);
	t(33) := t(10) - t(2);
	t(2) := fix_mul(924731744, t(33)) * 2;
	t(10) := t(11) + t(3);
	t(33) := t(11) - t(3);
	t(3) := fix_mul(684664577, t(33)) * 8;
	t(11) := t(12) + t(4);
	t(33) := t(12) - t(4);
	t(4) := fix_mul(608751522, t(33));
	t(12) := t(13) + t(5);
	t(33) := t(13) - t(5);
	t(5) := fix_mul(694519601, t(33));
	t(13) := t(14) + t(6);
	t(33) := t(14) - t(6);
	t(6) := fix_mul(561028615, t(33));
	t(14) := t(15) + t(7);
	t(33) := t(15) - t(7);
	t(7) := fix_mul(539468600, t(33));
	t(15) := t(4) + t(0);
	t(33) := t(4) - t(0);
	t(0) := fix_mul(966342111, t(33));
	t(4) := t(5) + t(1);
	t(33) := t(5) - t(1);
	t(1) := fix_mul(687977376, t(33)) * 4;
	t(5) := t(6) + t(2);
	t(33) := t(6) - t(2);
	t(2) := fix_mul(645689155, t(33));
	t(6) := t(7) + t(3);
	t(33) := t(7) - t(3);
	t(3) := fix_mul(547388834, t(33));
	t(7) := t(2) + t(0);
	t(33) := t(2) - t(0);
	t(0) := fix_mul(701455650, t(33)) * 2;
	t(2) := t(3) + t(1);
	t(33) := t(3) - t(1);
	t(1) := fix_mul(581104887, t(33));
	t(3) := t(1) + t(0);
	t(33) := t(1) - t(0);
	t(0) := fix_mul(759250124, t(33));
	t(1) := t(2) + t(7);
	t(33) := t(2) - t(7);
	t(2) := fix_mul(759250124, t(33));
	t(7) := t(0);
	t(3) := t(3) + t(0);
	t(0) := t(5) + t(15);
	t(33) := t(5) - t(15);
	t(5) := fix_mul(701455650, t(33)) * 2;
	t(15) := t(6) + t(4);
	t(33) := t(6) - t(4);
	t(4) := fix_mul(581104887, t(33));
	t(6) := t(4) + t(5);
	t(33) := t(4) - t(5);
	t(4) := fix_mul(759250124, t(33));
	t(5) := t(15) + t(0);
	t(33) := t(15) - t(0);
	t(0) := fix_mul(759250124, t(33));
	t(15) := t(4);
	t(6) := t(6) + t(4);
	t(4) := t(7);
	t(33) := t(7);
	t(7) := t(3);
	t(1) := t(1) + t(3);
	t(33) := t(33) + t(2);
	t(7) := t(7) + t(2);
	t(2) := t(11) + t(31);
	t(3) := t(11) - t(31);
	t(11) := fix_mul(966342111, t(3));
	t(3) := t(12) + t(8);
	t(31) := t(12) - t(8);
	t(8) := fix_mul(687977376, t(31)) * 4;
	t(12) := t(13) + t(9);
	t(31) := t(13) - t(9);
	t(9) := fix_mul(645689155, t(31));
	t(13) := t(14) + t(10);
	t(31) := t(14) - t(10);
	t(10) := fix_mul(547388834, t(31));
	t(14) := t(9) + t(11);
	t(31) := t(9) - t(11);
	t(9) := fix_mul(701455650, t(31)) * 2;
	t(11) := t(10) + t(8);
	t(31) := t(10) - t(8);
	t(8) := fix_mul(581104887, t(31));
	t(10) := t(8) + t(9);
	t(31) := t(8) - t(9);
	t(8) := fix_mul(759250124, t(31));
	t(9) := t(11) + t(14);
	t(31) := t(11) - t(14);
	t(11) := fix_mul(759250124, t(31));
	t(14) := t(8);
	t(10) := t(10) + t(8);
	t(8) := t(12) + t(2);
	t(31) := t(12) - t(2);
	t(2) := fix_mul(701455650, t(31)) * 2;
	t(12) := t(13) + t(3);
	t(31) := t(13) - t(3);
	t(3) := fix_mul(581104887, t(31));
	t(13) := t(3) + t(2);
	t(31) := t(3) - t(2);
	t(2) := fix_mul(759250124, t(31));
	t(3) := t(12) + t(8);
	t(31) := t(12) - t(8);
	t(8) := fix_mul(759250124, t(31));
	t(12) := t(2);
	t(13) := t(13) + t(2);
	t(2) := t(14);
	t(31) := t(14);
	t(14) := t(10);
	t(9) := t(9) + t(10);
	t(31) := t(31) + t(11);
	t(14) := t(14) + t(11);
	t(10) := t(4);
	t(11) := t(4);
	t(4) := t(7);
	t(34) := t(7);
	t(7) := t(33);
	t(35) := t(33);
	t(33) := t(1);
	t(5) := t(5) + t(1);
	t(11) := t(11) + t(15);
	t(7) := t(7) + t(15);
	t(34) := t(34) + t(6);
	t(33) := t(33) + t(6);
	t(35) := t(35) + t(0);
	t(4) := t(4) + t(0);
	t(0) := t(23) + t(32);
	t(1) := t(23) - t(32);
	t(6) := fix_mul(569446996, t(1)) * 2;
	t(1) := t(24) + t(16);
	t(15) := t(24) - t(16);
	t(16) := fix_mul(846274582, t(15));
	t(15) := t(25) + t(17);
	t(23) := t(25) - t(17);
	t(17) := fix_mul(924731744, t(23)) * 2;
	t(23) := t(26) + t(18);
	t(24) := t(26) - t(18);
	t(18) := fix_mul(684664577, t(24)) * 8;
	t(24) := t(27) + t(19);
	t(25) := t(27) - t(19);
	t(19) := fix_mul(608751522, t(25));
	t(25) := t(28) + t(20);
	t(26) := t(28) - t(20);
	t(20) := fix_mul(694519601, t(26));
	t(26) := t(29) + t(21);
	t(27) := t(29) - t(21);
	t(21) := fix_mul(561028615, t(27));
	t(27) := t(30) + t(22);
	t(28) := t(30) - t(22);
	t(22) := fix_mul(539468600, t(28));
	t(28) := t(19) + t(6);
	t(29) := t(19) - t(6);
	t(6) := fix_mul(966342111, t(29));
	t(19) := t(20) + t(16);
	t(29) := t(20) - t(16);
	t(16) := fix_mul(687977376, t(29)) * 4;
	t(20) := t(21) + t(17);
	t(29) := t(21) - t(17);
	t(17) := fix_mul(645689155, t(29));
	t(21) := t(22) + t(18);
	t(29) := t(22) - t(18);
	t(18) := fix_mul(547388834, t(29));
	t(22) := t(17) + t(6);
	t(29) := t(17) - t(6);
	t(6) := fix_mul(701455650, t(29)) * 2;
	t(17) := t(18) + t(16);
	t(29) := t(18) - t(16);
	t(16) := fix_mul(581104887, t(29));
	t(18) := t(16) + t(6);
	t(29) := t(16) - t(6);
	t(6) := fix_mul(759250124, t(29));
	t(16) := t(17) + t(22);
	t(29) := t(17) - t(22);
	t(17) := fix_mul(759250124, t(29));
	t(22) := t(6);
	t(18) := t(18) + t(6);
	t(6) := t(20) + t(28);
	t(29) := t(20) - t(28);
	t(20) := fix_mul(701455650, t(29)) * 2;
	t(28) := t(21) + t(19);
	t(29) := t(21) - t(19);
	t(19) := fix_mul(581104887, t(29));
	t(21) := t(19) + t(20);
	t(29) := t(19) - t(20);
	t(19) := fix_mul(759250124, t(29));
	t(20) := t(28) + t(6);
	t(29) := t(28) - t(6);
	t(6) := fix_mul(759250124, t(29));
	t(28) := t(19);
	t(21) := t(21) + t(19);
	t(19) := t(22);
	t(29) := t(22);
	t(22) := t(18);
	t(16) := t(16) + t(18);
	t(29) := t(29) + t(17);
	t(22) := t(22) + t(17);
	t(17) := t(24) + t(0);
	t(18) := t(24) - t(0);
	t(0) := fix_mul(966342111, t(18));
	t(18) := t(25) + t(1);
	t(24) := t(25) - t(1);
	t(1) := fix_mul(687977376, t(24)) * 4;
	t(24) := t(26) + t(15);
	t(25) := t(26) - t(15);
	t(15) := fix_mul(645689155, t(25));
	t(25) := t(27) + t(23);
	t(26) := t(27) - t(23);
	t(23) := fix_mul(547388834, t(26));
	t(26) := t(15) + t(0);
	t(27) := t(15) - t(0);
	t(0) := fix_mul(701455650, t(27)) * 2;
	t(15) := t(23) + t(1);
	t(27) := t(23) - t(1);
	t(1) := fix_mul(581104887, t(27));
	t(23) := t(1) + t(0);
	t(27) := t(1) - t(0);
	t(0) := fix_mul(759250124, t(27));
	t(1) := t(15) + t(26);
	t(27) := t(15) - t(26);
	t(15) := fix_mul(759250124, t(27));
	t(26) := t(0);
	t(23) := t(23) + t(0);
	t(0) := t(24) + t(17);
	t(27) := t(24) - t(17);
	t(17) := fix_mul(701455650, t(27)) * 2;
	t(24) := t(25) + t(18);
	t(27) := t(25) - t(18);
	t(18) := fix_mul(581104887, t(27));
	t(25) := t(18) + t(17);
	t(27) := t(18) - t(17);
	t(17) := fix_mul(759250124, t(27));
	t(18) := t(24) + t(0);
	t(27) := t(24) - t(0);
	t(0) := fix_mul(759250124, t(27));
	t(24) := t(17);
	t(25) := t(25) + t(17);
	t(17) := t(26);
	t(27) := t(26);
	t(26) := t(23);
	t(1) := t(1) + t(23);
	t(27) := t(27) + t(15);
	t(26) := t(26) + t(15);
	t(15) := t(19);
	t(23) := t(19);
	t(19) := t(22);
	t(30) := t(22);
	t(22) := t(29);
	t(32) := t(29);
	t(29) := t(16);
	t(20) := t(20) + t(16);
	t(23) := t(23) + t(28);
	t(22) := t(22) + t(28);
	t(30) := t(30) + t(21);
	t(29) := t(29) + t(21);
	t(32) := t(32) + t(6);
	t(19) := t(19) + t(6);
	t(6) := t(10);
	t(16) := t(10);
	t(10) := t(4);
	t(21) := t(4);
	t(4) := t(7);
	t(28) := t(7);
	t(7) := t(33);
	t(36) := t(33);
	t(33) := t(11);
	t(37) := t(11);
	t(11) := t(34);
	t(38) := t(34);
	t(34) := t(35);
	t(39) := t(35);
	t(35) := t(5);
	t(3) := t(3) + t(5);
	t(16) := t(16) + t(2);
	t(33) := t(33) + t(2);
	t(21) := t(21) + t(14);
	t(11) := t(11) + t(14);
	t(28) := t(28) + t(31);
	t(34) := t(34) + t(31);
	t(36) := t(36) + t(9);
	t(35) := t(35) + t(9);
	t(37) := t(37) + t(12);
	t(4) := t(4) + t(12);
	t(38) := t(38) + t(13);
	t(7) := t(7) + t(13);
	t(39) := t(39) + t(8);
	t(10) := t(10) + t(8);
	VOffsetPtr(0) := 0-t(6);
	VOffsetPtr(1) := 0-t(10);
	VOffsetPtr(2) := 0-t(4);
	VOffsetPtr(3) := 0-t(7);
	VOffsetPtr(4) := 0-t(33);
	VOffsetPtr(5) := 0-t(11);
	VOffsetPtr(6) := 0-t(34);
	VOffsetPtr(7) := 0-t(35);
	VOffsetPtr(8) := 0-t(16);
	VOffsetPtr(9) := 0-t(21);
	VOffsetPtr(10) := 0-t(28);
	VOffsetPtr(11) := 0-t(36);
	VOffsetPtr(12) := 0-t(37);
	VOffsetPtr(13) := 0-t(38);
	VOffsetPtr(14) := 0-t(39);
	VOffsetPtr(15) := 0-t(3);
	VOffsetPtr(16) := 0-t(15);
	VOffsetPtr(17) := 0-t(19);
	VOffsetPtr(18) := 0-t(22);
	VOffsetPtr(19) := 0-t(29);
	VOffsetPtr(20) := 0-t(23);
	VOffsetPtr(21) := 0-t(30);
	VOffsetPtr(22) := 0-t(32);
	VOffsetPtr(23) := 0-t(20);
	VOffsetPtr(24) := 0-t(17);
	VOffsetPtr(25) := 0-t(26);
	VOffsetPtr(26) := 0-t(27);
	VOffsetPtr(27) := 0-t(1);
	VOffsetPtr(28) := 0-t(24);
	VOffsetPtr(29) := 0-t(25);
	VOffsetPtr(30) := 0-t(0);
	VOffsetPtr(31) := 0-t(18);
	
	return VOffsetPtr;
     end;
	
end;
�