-- 
-- psg_wave.vhd
--   Programmable Sound Generator (AY-3-8910/YM2149)
--   Revision 1.00
-- 
-- Copyright (c) 2006 Kazuhiro Tsujikawa (ESE Artists' factory)
-- All rights reserved.
-- 
-- Redistribution and use of this source code or any derivative works, are 
-- permitted provided that the following conditions are met:
--
-- 1. Redistributions of source code must retain the above copyright notice, 
--    this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright 
--    notice, this list of conditions and the following disclaimer in the 
--    documentation and/or other materials provided with the distribution.
-- 3. Redistributions may not be sold, nor may they be used in a commercial 
--    product or activity without specific prior written permission.
--
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS 
-- "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED 
-- TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR 
-- PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT OWNER OR 
-- CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, 
-- EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, 
-- PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS;
-- OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, 
-- WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR 
-- OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF 
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 

LIBRARY IEEE;
	USE IEEE.STD_LOGIC_1164.ALL;
	USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PSG_WAVE IS
	PORT(
		CLK21M		: IN	STD_LOGIC;
		RESET		: IN	STD_LOGIC;
		CLKENA		: IN	STD_LOGIC;
		REQ			: IN	STD_LOGIC;
		ACK			: OUT	STD_LOGIC;
		WRT			: IN	STD_LOGIC;
		ADR			: IN	STD_LOGIC_VECTOR( 15 DOWNTO 0 );
		DBI			: OUT	STD_LOGIC_VECTOR(  7 DOWNTO 0 );
		DBO			: IN	STD_LOGIC_VECTOR(  7 DOWNTO 0 );
		WAVE		: OUT	STD_LOGIC_VECTOR(  7 DOWNTO 0 )
	);
END PSG_WAVE;

ARCHITECTURE RTL OF PSG_WAVE IS

	SIGNAL PSGCLKENA	: STD_LOGIC_VECTOR(  4 DOWNTO 0 );
	SIGNAL PSGREGPTR	: STD_LOGIC_VECTOR(  3 DOWNTO 0 );

	SIGNAL PSGEDGECHA	: STD_LOGIC;
	SIGNAL PSGEDGECHB	: STD_LOGIC;
	SIGNAL PSGEDGECHC	: STD_LOGIC;
	SIGNAL PSGNOISE		: STD_LOGIC;
	SIGNAL PSGVOLENV	: STD_LOGIC_VECTOR(  3 DOWNTO 0 );
	SIGNAL PSGENVREQ	: STD_LOGIC;
	SIGNAL PSGENVACK	: STD_LOGIC;

	SIGNAL PSGFREQCHA	: STD_LOGIC_VECTOR( 11 DOWNTO 0 );
	SIGNAL PSGFREQCHB	: STD_LOGIC_VECTOR( 11 DOWNTO 0 );
	SIGNAL PSGFREQCHC	: STD_LOGIC_VECTOR( 11 DOWNTO 0 );
	SIGNAL PSGFREQNOISE	: STD_LOGIC_VECTOR(  4 DOWNTO 0 );
	SIGNAL PSGCHANSEL	: STD_LOGIC_VECTOR(  5 DOWNTO 0 );
	SIGNAL PSGVOLCHA	: STD_LOGIC_VECTOR(  4 DOWNTO 0 );
	SIGNAL PSGVOLCHB	: STD_LOGIC_VECTOR(  4 DOWNTO 0 );
	SIGNAL PSGVOLCHC	: STD_LOGIC_VECTOR(  4 DOWNTO 0 );
	SIGNAL PSGFREQENV	: STD_LOGIC_VECTOR( 15 DOWNTO 0 );
	SIGNAL PSGSHAPEENV	: STD_LOGIC_VECTOR(  3 DOWNTO 0 );

	ALIAS HOLD			: STD_LOGIC IS PSGSHAPEENV(0);
	ALIAS ALTER			: STD_LOGIC IS PSGSHAPEENV(1);
	ALIAS ATTACK		: STD_LOGIC IS PSGSHAPEENV(2);
	ALIAS CONT			: STD_LOGIC IS PSGSHAPEENV(3);

BEGIN

	----------------------------------------------------------------
	-- MISCELLANEOUS CONTROL / CLOCK ENABLE (DIVIDER)
	----------------------------------------------------------------
	PROCESS( RESET, CLK21M )
	BEGIN
		IF( RESET = '1' )THEN
			PSGCLKENA <= (OTHERS => '0');
		ELSIF (CLK21M'EVENT AND CLK21M = '1') THEN
			IF( CLKENA = '1' )THEN
				PSGCLKENA <= PSGCLKENA - 1;
			END IF;
		END IF;
	END PROCESS;

	ACK <= REQ;

	----------------------------------------------------------------
	-- PSG REGISTER READ
	----------------------------------------------------------------
	DBI <=					PSGFREQCHA( 7 DOWNTO 0) WHEN( PSGREGPTR = "0000" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"0000"	&	PSGFREQCHA(11 DOWNTO 8) WHEN( PSGREGPTR = "0001" AND ADR(1 DOWNTO 0) = "10" )ELSE
							PSGFREQCHB( 7 DOWNTO 0) WHEN( PSGREGPTR = "0010" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"0000"	&	PSGFREQCHB(11 DOWNTO 8) WHEN( PSGREGPTR = "0011" AND ADR(1 DOWNTO 0) = "10" )ELSE
							PSGFREQCHC( 7 DOWNTO 0) WHEN( PSGREGPTR = "0100" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"0000"	&	PSGFREQCHC(11 DOWNTO 8) WHEN( PSGREGPTR = "0101" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"000"	&	PSGFREQNOISE			WHEN( PSGREGPTR = "0110" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"10"	&	PSGCHANSEL				WHEN( PSGREGPTR = "0111" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"000"	&	PSGVOLCHA				WHEN( PSGREGPTR = "1000" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"000"	&	PSGVOLCHB				WHEN( PSGREGPTR = "1001" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"000"	&	PSGVOLCHC				WHEN( PSGREGPTR = "1010" AND ADR(1 DOWNTO 0) = "10" )ELSE
				PSGFREQENV(7 DOWNTO 0)				WHEN( PSGREGPTR = "1011" AND ADR(1 DOWNTO 0) = "10" )ELSE
				PSGFREQENV(15 DOWNTO 8)				WHEN( PSGREGPTR = "1100" AND ADR(1 DOWNTO 0) = "10" )ELSE
				"0000" & PSGSHAPEENV				WHEN( PSGREGPTR = "1101" AND ADR(1 DOWNTO 0) = "10" )ELSE
				(OTHERS => '1');

	----------------------------------------------------------------
	-- PSG REGISTER WRITE
	----------------------------------------------------------------
	PROCESS(CLK21M, RESET)

	BEGIN

		IF (RESET = '1') THEN

			PSGREGPTR		 <= (OTHERS => '0');

			PSGFREQCHA	 <= (OTHERS => '1');
			PSGFREQCHB	 <= (OTHERS => '1');
			PSGFREQCHC	 <= (OTHERS => '1');
			PSGFREQNOISE <= (OTHERS => '1');
			PSGCHANSEL	 <= (OTHERS => '1');
			PSGVOLCHA		 <= (OTHERS => '1');
			PSGVOLCHB		 <= (OTHERS => '1');
			PSGVOLCHC		 <= (OTHERS => '1');
			PSGFREQENV	 <= (OTHERS => '1');
			PSGSHAPEENV	 <= (OTHERS => '1');
			PSGENVREQ		 <= '0';

		ELSIF (CLK21M'EVENT AND CLK21M = '1') THEN

			IF (REQ = '1' AND WRT = '1' AND ADR(1 DOWNTO 0) = "00") THEN
				-- REGISTER POINTER
				PSGREGPTR <= DBO(3 DOWNTO 0);
			ELSIF (REQ = '1' AND WRT = '1' AND ADR(1 DOWNTO 0) = "01") THEN
				-- PSG REGISTERS
				CASE PSGREGPTR IS
					WHEN "0000" => PSGFREQCHA(7 DOWNTO 0)	 <= DBO;
					WHEN "0001" => PSGFREQCHA(11 DOWNTO 8) <= DBO(3 DOWNTO 0);
					WHEN "0010" => PSGFREQCHB(7 DOWNTO 0)	 <= DBO;
					WHEN "0011" => PSGFREQCHB(11 DOWNTO 8) <= DBO(3 DOWNTO 0);
					WHEN "0100" => PSGFREQCHC(7 DOWNTO 0)	 <= DBO;
					WHEN "0101" => PSGFREQCHC(11 DOWNTO 8) <= DBO(3 DOWNTO 0);
					WHEN "0110" => PSGFREQNOISE						 <= DBO(4 DOWNTO 0);
					WHEN "0111" => PSGCHANSEL							 <= DBO(5 DOWNTO 0);
					WHEN "1000" => PSGVOLCHA							 <= DBO(4 DOWNTO 0);
					WHEN "1001" => PSGVOLCHB							 <= DBO(4 DOWNTO 0);
					WHEN "1010" => PSGVOLCHC							 <= DBO(4 DOWNTO 0);
					WHEN "1011" => PSGFREQENV(7 DOWNTO 0)	 <= DBO;
					WHEN "1100" => PSGFREQENV(15 DOWNTO 8) <= DBO;
					WHEN "1101" => PSGSHAPEENV						 <= DBO(3 DOWNTO 0); PSGENVREQ <= NOT PSGENVACK;
					WHEN OTHERS => NULL;
				END CASE;
			END IF;

		END IF;

	END PROCESS;

	----------------------------------------------------------------
	-- TONE GENERATOR
	----------------------------------------------------------------
	PROCESS(CLK21M, RESET)

		VARIABLE PSGCNTCHA : STD_LOGIC_VECTOR(11 DOWNTO 0);
		VARIABLE PSGCNTCHB : STD_LOGIC_VECTOR(11 DOWNTO 0);
		VARIABLE PSGCNTCHC : STD_LOGIC_VECTOR(11 DOWNTO 0);

	BEGIN

		IF (RESET = '1') THEN

			PSGEDGECHA <= '0';
			PSGCNTCHA	 := (OTHERS => '0');
			PSGEDGECHB <= '0';
			PSGCNTCHB	 := (OTHERS => '0');
			PSGEDGECHC <= '0';
			PSGCNTCHC	 := (OTHERS => '0');

		ELSIF (CLK21M'EVENT AND CLK21M = '1') THEN

			-- BASE FREQUENCY : 112KHZ = 3.58MHZ / 16 / 2
			IF (PSGCLKENA(3 DOWNTO 0) = "0000" AND CLKENA = '1') THEN

				IF (PSGCNTCHA /= X"000") THEN
					PSGCNTCHA := PSGCNTCHA - 1;
				ELSIF (PSGFREQCHA /= X"000") THEN
					PSGCNTCHA := PSGFREQCHA - 1;
				END IF;
				IF (PSGCNTCHA = X"000") THEN
					PSGEDGECHA <= NOT PSGEDGECHA;
				END IF;

				IF (PSGCNTCHB /= X"000") THEN
					PSGCNTCHB := PSGCNTCHB - 1;
				ELSIF (PSGFREQCHB /= X"000") THEN
					PSGCNTCHB := PSGFREQCHB - 1;
				END IF;
				IF (PSGCNTCHB = X"000") THEN
					PSGEDGECHB <= NOT PSGEDGECHB;
				END IF;

				IF (PSGCNTCHC /= X"000") THEN
					PSGCNTCHC := PSGCNTCHC - 1;
				ELSIF (PSGFREQCHC /= X"000") THEN
					PSGCNTCHC := PSGFREQCHC - 1;
				END IF;
				IF (PSGCNTCHC = X"000") THEN
					PSGEDGECHC <= NOT PSGEDGECHC;
				END IF;

			END IF;

		END IF;

	END PROCESS;

	----------------------------------------------------------------
	-- NOISE GENERATOR 
	----------------------------------------------------------------
	PROCESS(CLK21M, RESET)

		VARIABLE PSGCNTNOISE : STD_LOGIC_VECTOR(4 DOWNTO 0);
		VARIABLE PSGGENNOISE : STD_LOGIC_VECTOR(17 DOWNTO 0);

	BEGIN

		IF (RESET = '1') THEN

			PSGCNTNOISE := (OTHERS => '0');
			PSGGENNOISE := (OTHERS => '1');

		ELSIF (CLK21M'EVENT AND CLK21M = '1') THEN

			-- BASE FREQUENCY : 112KHZ = 3.58MHZ / 16 / 2
			IF (PSGCLKENA(4 DOWNTO 0) = "00000" AND CLKENA = '1') THEN

				-- NOISE FREQUENCY COUNTER
				IF (PSGCNTNOISE /= "00000") THEN
					PSGCNTNOISE := PSGCNTNOISE - 1;
				ELSIF (PSGFREQNOISE /= "00000") THEN
					PSGCNTNOISE := PSGFREQNOISE - 1;
				END IF;

				-- (MAXIMUM-LENGTH LINEAR SHIFT REGISTER SEQUENCE)
				-- F(X) = X^17 + X^14 + 1
				IF (PSGCNTNOISE = "00000") THEN

					FOR I IN 17 DOWNTO 1 LOOP
						PSGGENNOISE(I) := PSGGENNOISE(I - 1);
					END LOOP;

					IF (PSGGENNOISE = "00000000000000000") THEN
						PSGGENNOISE(0) := '1';																					-- ERROR TRAP
					ELSE
						PSGGENNOISE(0) := PSGGENNOISE(17) XOR PSGGENNOISE(14);					-- NORMAL WORK
					END IF;

				END IF;

			END IF;

		END IF;

		PSGNOISE <= PSGGENNOISE(17);

	END PROCESS;

	----------------------------------------------------------------
	-- ENVELOPE GENERATOR
	----------------------------------------------------------------
	PROCESS(CLK21M, RESET)

		VARIABLE PSGCNTENV : STD_LOGIC_VECTOR(15 DOWNTO 0);
		VARIABLE PSGPTRENV : STD_LOGIC_VECTOR(4 DOWNTO 0);

	BEGIN

		IF (RESET = '1') THEN

			PSGCNTENV := (OTHERS => '0');
			PSGPTRENV := (OTHERS => '1');
			PSGVOLENV <= (OTHERS => '0');
			PSGENVACK <= '0';

		ELSIF (CLK21M'EVENT AND CLK21M = '1') THEN

			-- ENVELOPE BASE FREQUENCY : 56KHZ = 3.58MHZ / 8 / 2
			IF (PSGCLKENA(4 DOWNTO 0) = "00000" AND CLKENA = '1') THEN

				-- ENVELOPE PREIOD COUNTER
				IF (PSGCNTENV /= X"0000" AND PSGENVREQ = PSGENVACK) THEN
					PSGCNTENV := PSGCNTENV - 1;
				ELSIF (PSGFREQENV /= X"0000") THEN
					PSGCNTENV := PSGFREQENV - 1;
				END IF;

				-- ENVELOPE PHASE COUNTER
				IF (PSGENVREQ /= PSGENVACK) THEN
					PSGPTRENV := (OTHERS => '1');
				ELSIF (PSGCNTENV = X"0000" AND (PSGPTRENV(4) = '1' OR (HOLD = '0' AND CONT = '1'))) THEN
					PSGPTRENV := PSGPTRENV - 1;
				END IF;

				-- ENVELOPE AMPLITUDE CONTROL
				FOR I IN 3 DOWNTO 0 LOOP
					IF (PSGPTRENV(4) = '0' AND CONT = '0') THEN
						PSGVOLENV(I) <= '0';
					ELSIF (PSGPTRENV(4) = '1' OR (ALTER XOR HOLD) = '0') THEN
						PSGVOLENV(I) <= PSGPTRENV(I) XOR ATTACK;
					ELSE
						PSGVOLENV(I) <= PSGPTRENV(I) XOR ATTACK XOR '1';
					END IF;
				END LOOP;

				PSGENVACK <= PSGENVREQ;

			END IF;

		END IF;

	END PROCESS;

	----------------------------------------------------------------
	-- MIXER CONTROL
	----------------------------------------------------------------
	PROCESS(CLK21M, RESET)

		VARIABLE PSGENANOISE : STD_LOGIC;
		VARIABLE PSGENATONE	 : STD_LOGIC;
		VARIABLE PSGEDGE		 : STD_LOGIC;
		VARIABLE PSGVOL			 : STD_LOGIC_VECTOR(4 DOWNTO 0);
		VARIABLE PSGINDEX		 : STD_LOGIC_VECTOR(3 DOWNTO 0);
		VARIABLE PSGTABLE		 : STD_LOGIC_VECTOR(7 DOWNTO 0);
		VARIABLE PSGMIX			 : STD_LOGIC_VECTOR(9 DOWNTO 0);

	BEGIN

		IF (RESET = '1') THEN

			PSGMIX := (OTHERS => '0');
			WAVE	 <= (OTHERS => '0');

		ELSIF (CLK21M'EVENT AND CLK21M = '1') THEN

			CASE PSGCLKENA(1 DOWNTO 0) IS
				WHEN "11"		=>
					PSGENATONE	:= PSGCHANSEL(0); PSGEDGE	 := PSGEDGECHA;
					PSGENANOISE := PSGCHANSEL(3); PSGVOL	 := PSGVOLCHA;
				WHEN "10"		=>
					PSGENATONE	:= PSGCHANSEL(1); PSGEDGE	 := PSGEDGECHB;
					PSGENANOISE := PSGCHANSEL(4); PSGVOL	 := PSGVOLCHB;
				WHEN "01"		=>
					PSGENATONE	:= PSGCHANSEL(2); PSGEDGE	 := PSGEDGECHC;
					PSGENANOISE := PSGCHANSEL(5); PSGVOL	 := PSGVOLCHC;
				WHEN OTHERS =>
					PSGENATONE	:= '1';						PSGEDGE	 := '1';
					PSGENANOISE := '1';						PSGVOL	 := "00000";
			END CASE;

			IF (((PSGENATONE OR PSGEDGE) AND (PSGENANOISE OR PSGNOISE)) = '0') THEN
				PSGINDEX := (OTHERS => '0');
			ELSIF (PSGVOL(4) = '0') THEN
				PSGINDEX := PSGVOL(3 DOWNTO 0);
			ELSE
				PSGINDEX := PSGVOLENV;
			END IF;

			CASE PSGINDEX IS
				WHEN "1111" => PSGTABLE := "11111111";
				WHEN "1110" => PSGTABLE := "10110100";
				WHEN "1101" => PSGTABLE := "01111111";
				WHEN "1100" => PSGTABLE := "01011010";
				WHEN "1011" => PSGTABLE := "00111111";
				WHEN "1010" => PSGTABLE := "00101101";
				WHEN "1001" => PSGTABLE := "00011111";
				WHEN "1000" => PSGTABLE := "00010110";
				WHEN "0111" => PSGTABLE := "00001111";
				WHEN "0110" => PSGTABLE := "00001011";
				WHEN "0101" => PSGTABLE := "00000111";
				WHEN "0100" => PSGTABLE := "00000101";
				WHEN "0011" => PSGTABLE := "00000011";
				WHEN "0010" => PSGTABLE := "00000010";
				WHEN "0001" => PSGTABLE := "00000001";
				WHEN OTHERS => PSGTABLE := "00000000";
			END CASE;

			IF (CLKENA = '1') THEN
				CASE PSGCLKENA(1 DOWNTO 0) IS
					WHEN "00"		=> WAVE		<= PSGMIX(9 DOWNTO 2);
												 PSGMIX(9 DOWNTO 2) := (OTHERS => '0');
					WHEN OTHERS => PSGMIX := "00" & PSGTABLE + PSGMIX;
				END CASE;
			END IF;

		END IF;

	END PROCESS;

END RTL;
