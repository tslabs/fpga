`timescale 1ns / 1ps

module ssram(
	input	wire		CLK,
	
	input	wire [14:0]	ADDR, //16kb
	input	wire [7:0]	DI,
	output	wire [7:0]	DO,
	input	wire		OE,
	input	wire		WE
); 	   

reg [7:0]	ram [0:32*1024-1];

always @ (negedge CLK)
if (WE)		 	
begin
	ram[ADDR] = DI;
	//$display("MEM WRITE ADDR=%h VAL=%h", ADDR, DI);
end
	
assign #1 DO = ram[ADDR];

integer i;

initial
begin	
		for(i=0;i<32*1024;i=i+1)
			ram[i] = 0;
	

		
		ram[15'h0] =  8'hC3;
		ram[15'h1] =  8'h4B;
		ram[15'h2] =  8'h00;
		ram[15'h3] =  8'h00;
		ram[15'h4] =  8'h00;
		ram[15'h5] =  8'h00;
		ram[15'h6] =  8'h00;
		ram[15'h7] =  8'h00;
		ram[15'h8] =  8'h00;
		ram[15'h9] =  8'h00;
		ram[15'hA] =  8'h00;
		ram[15'hB] =  8'h00;
		ram[15'hC] =  8'h00;
		ram[15'hD] =  8'h00;
		ram[15'hE] =  8'h00;
		ram[15'hF] =  8'h00;
		ram[15'h10] =  8'hD3;
		ram[15'h11] =  8'hFF;
		ram[15'h12] =  8'hC9;
		ram[15'h13] =  8'h00;
		ram[15'h14] =  8'h00;
		ram[15'h15] =  8'h00;
		ram[15'h16] =  8'h00;
		ram[15'h17] =  8'h00;
		ram[15'h18] =  8'h00;
		ram[15'h19] =  8'h00;
		ram[15'h1A] =  8'h00;
		ram[15'h1B] =  8'h00;
		ram[15'h1C] =  8'h00;
		ram[15'h1D] =  8'h00;
		ram[15'h1E] =  8'h00;
		ram[15'h1F] =  8'h00;
		ram[15'h20] =  8'h00;
		ram[15'h21] =  8'h00;
		ram[15'h22] =  8'h00;
		ram[15'h23] =  8'h00;
		ram[15'h24] =  8'h00;
		ram[15'h25] =  8'h00;
		ram[15'h26] =  8'h00;
		ram[15'h27] =  8'h00;
		ram[15'h28] =  8'h00;
		ram[15'h29] =  8'h00;
		ram[15'h2A] =  8'h00;
		ram[15'h2B] =  8'h00;
		ram[15'h2C] =  8'h00;
		ram[15'h2D] =  8'h00;
		ram[15'h2E] =  8'h00;
		ram[15'h2F] =  8'h00;
		ram[15'h30] =  8'h00;
		ram[15'h31] =  8'h00;
		ram[15'h32] =  8'h00;
		ram[15'h33] =  8'h00;
		ram[15'h34] =  8'h00;
		ram[15'h35] =  8'h00;
		ram[15'h36] =  8'h00;
		ram[15'h37] =  8'h00;
		ram[15'h38] =  8'hED;
		ram[15'h39] =  8'h4D;
		ram[15'h3A] =  8'h00;
		ram[15'h3B] =  8'h00;
		ram[15'h3C] =  8'h00;
		ram[15'h3D] =  8'h00;
		ram[15'h3E] =  8'h00;
		ram[15'h3F] =  8'h00;
		ram[15'h40] =  8'h00;
		ram[15'h41] =  8'h00;
		ram[15'h42] =  8'h00;
		ram[15'h43] =  8'h00;
		ram[15'h44] =  8'h00;
		ram[15'h45] =  8'h00;
		ram[15'h46] =  8'h00;
		ram[15'h47] =  8'h00;
		ram[15'h48] =  8'h00;
		ram[15'h49] =  8'h00;
		ram[15'h4A] =  8'hF5;
		ram[15'h4B] =  8'h21;
		ram[15'h4C] =  8'hFF;
		ram[15'h4D] =  8'h23;
		ram[15'h4E] =  8'hF9;
		ram[15'h4F] =  8'h11;
		ram[15'h50] =  8'h34;
		ram[15'h51] =  8'h1D;
		ram[15'h52] =  8'h0E;
		ram[15'h53] =  8'h09;
		ram[15'h54] =  8'hCD;
		ram[15'h55] =  8'h0C;
		ram[15'h56] =  8'h1D;
		ram[15'h57] =  8'h21;
		ram[15'h58] =  8'h72;
		ram[15'h59] =  8'h00;
		ram[15'h5A] =  8'h7E;
		ram[15'h5B] =  8'h23;
		ram[15'h5C] =  8'hB6;
		ram[15'h5D] =  8'hCA;
		ram[15'h5E] =  8'h67;
		ram[15'h5F] =  8'h00;
		ram[15'h60] =  8'h2B;
		ram[15'h61] =  8'hCD;
		ram[15'h62] =  8'h1A;
		ram[15'h63] =  8'h1A;
		ram[15'h64] =  8'hC3;
		ram[15'h65] =  8'h5A;
		ram[15'h66] =  8'h00;
		ram[15'h67] =  8'h11;
		ram[15'h68] =  8'h55;
		ram[15'h69] =  8'h1D;
		ram[15'h6A] =  8'h0E;
		ram[15'h6B] =  8'h09;
		ram[15'h6C] =  8'hCD;
		ram[15'h6D] =  8'h0C;
		ram[15'h6E] =  8'h1D;
		ram[15'h6F] =  8'hC3;
		ram[15'h70] =  8'h6F;
		ram[15'h71] =  8'h00;
		ram[15'h72] =  8'hFA;
		ram[15'h73] =  8'h00;
		ram[15'h74] =  8'h5A;
		ram[15'h75] =  8'h01;
		ram[15'h76] =  8'hBA;
		ram[15'h77] =  8'h01;
		ram[15'h78] =  8'h1A;
		ram[15'h79] =  8'h02;
		ram[15'h7A] =  8'h7A;
		ram[15'h7B] =  8'h02;
		ram[15'h7C] =  8'hDA;
		ram[15'h7D] =  8'h02;
		ram[15'h7E] =  8'h3A;
		ram[15'h7F] =  8'h03;
		ram[15'h80] =  8'h9A;
		ram[15'h81] =  8'h03;
		ram[15'h82] =  8'hFA;
		ram[15'h83] =  8'h03;
		ram[15'h84] =  8'h5A;
		ram[15'h85] =  8'h04;
		ram[15'h86] =  8'hBA;
		ram[15'h87] =  8'h04;
		ram[15'h88] =  8'h1A;
		ram[15'h89] =  8'h05;
		ram[15'h8A] =  8'h7A;
		ram[15'h8B] =  8'h05;
		ram[15'h8C] =  8'hDA;
		ram[15'h8D] =  8'h05;
		ram[15'h8E] =  8'h3A;
		ram[15'h8F] =  8'h06;
		ram[15'h90] =  8'h9A;
		ram[15'h91] =  8'h06;
		ram[15'h92] =  8'hFA;
		ram[15'h93] =  8'h06;
		ram[15'h94] =  8'h5A;
		ram[15'h95] =  8'h07;
		ram[15'h96] =  8'hBA;
		ram[15'h97] =  8'h07;
		ram[15'h98] =  8'h1A;
		ram[15'h99] =  8'h08;
		ram[15'h9A] =  8'h7A;
		ram[15'h9B] =  8'h08;
		ram[15'h9C] =  8'hDA;
		ram[15'h9D] =  8'h08;
		ram[15'h9E] =  8'h3A;
		ram[15'h9F] =  8'h09;
		ram[15'hA0] =  8'h9A;
		ram[15'hA1] =  8'h09;
		ram[15'hA2] =  8'hFA;
		ram[15'hA3] =  8'h09;
		ram[15'hA4] =  8'h5A;
		ram[15'hA5] =  8'h0A;
		ram[15'hA6] =  8'hBA;
		ram[15'hA7] =  8'h0A;
		ram[15'hA8] =  8'h1A;
		ram[15'hA9] =  8'h0B;
		ram[15'hAA] =  8'h7A;
		ram[15'hAB] =  8'h0B;
		ram[15'hAC] =  8'hDA;
		ram[15'hAD] =  8'h0B;
		ram[15'hAE] =  8'h3A;
		ram[15'hAF] =  8'h0C;
		ram[15'hB0] =  8'h9A;
		ram[15'hB1] =  8'h0C;
		ram[15'hB2] =  8'hFA;
		ram[15'hB3] =  8'h0C;
		ram[15'hB4] =  8'h5A;
		ram[15'hB5] =  8'h0D;
		ram[15'hB6] =  8'hBA;
		ram[15'hB7] =  8'h0D;
		ram[15'hB8] =  8'h1A;
		ram[15'hB9] =  8'h0E;
		ram[15'hBA] =  8'h7A;
		ram[15'hBB] =  8'h0E;
		ram[15'hBC] =  8'hDA;
		ram[15'hBD] =  8'h0E;
		ram[15'hBE] =  8'h3A;
		ram[15'hBF] =  8'h0F;
		ram[15'hC0] =  8'h9A;
		ram[15'hC1] =  8'h0F;
		ram[15'hC2] =  8'hFA;
		ram[15'hC3] =  8'h0F;
		ram[15'hC4] =  8'h5A;
		ram[15'hC5] =  8'h10;
		ram[15'hC6] =  8'hBA;
		ram[15'hC7] =  8'h10;
		ram[15'hC8] =  8'h1A;
		ram[15'hC9] =  8'h11;
		ram[15'hCA] =  8'h7A;
		ram[15'hCB] =  8'h11;
		ram[15'hCC] =  8'hDA;
		ram[15'hCD] =  8'h11;
		ram[15'hCE] =  8'h3A;
		ram[15'hCF] =  8'h12;
		ram[15'hD0] =  8'h9A;
		ram[15'hD1] =  8'h12;
		ram[15'hD2] =  8'hFA;
		ram[15'hD3] =  8'h12;
		ram[15'hD4] =  8'h5A;
		ram[15'hD5] =  8'h13;
		ram[15'hD6] =  8'hBA;
		ram[15'hD7] =  8'h13;
		ram[15'hD8] =  8'h1A;
		ram[15'hD9] =  8'h14;
		ram[15'hDA] =  8'h7A;
		ram[15'hDB] =  8'h14;
		ram[15'hDC] =  8'hDA;
		ram[15'hDD] =  8'h14;
		ram[15'hDE] =  8'h3A;
		ram[15'hDF] =  8'h15;
		ram[15'hE0] =  8'h9A;
		ram[15'hE1] =  8'h15;
		ram[15'hE2] =  8'hFA;
		ram[15'hE3] =  8'h15;
		ram[15'hE4] =  8'h5A;
		ram[15'hE5] =  8'h16;
		ram[15'hE6] =  8'hBA;
		ram[15'hE7] =  8'h16;
		ram[15'hE8] =  8'h1A;
		ram[15'hE9] =  8'h17;
		ram[15'hEA] =  8'h7A;
		ram[15'hEB] =  8'h17;
		ram[15'hEC] =  8'hDA;
		ram[15'hED] =  8'h17;
		ram[15'hEE] =  8'h3A;
		ram[15'hEF] =  8'h18;
		ram[15'hF0] =  8'h9A;
		ram[15'hF1] =  8'h18;
		ram[15'hF2] =  8'hFA;
		ram[15'hF3] =  8'h18;
		ram[15'hF4] =  8'h5A;
		ram[15'hF5] =  8'h19;
		ram[15'hF6] =  8'hBA;
		ram[15'hF7] =  8'h19;
		ram[15'hF8] =  8'h00;
		ram[15'hF9] =  8'h00;
		ram[15'hFA] =  8'hC7;
		ram[15'hFB] =  8'hED;
		ram[15'hFC] =  8'h42;
		ram[15'hFD] =  8'h00;
		ram[15'hFE] =  8'h00;
		ram[15'hFF] =  8'h2C;
		ram[15'h100] =  8'h83;
		ram[15'h101] =  8'h88;
		ram[15'h102] =  8'h4F;
		ram[15'h103] =  8'h2B;
		ram[15'h104] =  8'hF2;
		ram[15'h105] =  8'h39;
		ram[15'h106] =  8'hB3;
		ram[15'h107] =  8'h1F;
		ram[15'h108] =  8'h7E;
		ram[15'h109] =  8'h63;
		ram[15'h10A] =  8'h15;
		ram[15'h10B] =  8'hD3;
		ram[15'h10C] =  8'h89;
		ram[15'h10D] =  8'h5E;
		ram[15'h10E] =  8'h46;
		ram[15'h10F] =  8'h00;
		ram[15'h110] =  8'h38;
		ram[15'h111] =  8'h00;
		ram[15'h112] =  8'h00;
		ram[15'h113] =  8'h00;
		ram[15'h114] =  8'h00;
		ram[15'h115] =  8'h00;
		ram[15'h116] =  8'h00;
		ram[15'h117] =  8'h00;
		ram[15'h118] =  8'h00;
		ram[15'h119] =  8'h21;
		ram[15'h11A] =  8'hF8;
		ram[15'h11B] =  8'h00;
		ram[15'h11C] =  8'h00;
		ram[15'h11D] =  8'h00;
		ram[15'h11E] =  8'h00;
		ram[15'h11F] =  8'h00;
		ram[15'h120] =  8'h00;
		ram[15'h121] =  8'h00;
		ram[15'h122] =  8'h00;
		ram[15'h123] =  8'h00;
		ram[15'h124] =  8'h00;
		ram[15'h125] =  8'h00;
		ram[15'h126] =  8'h00;
		ram[15'h127] =  8'h00;
		ram[15'h128] =  8'h00;
		ram[15'h129] =  8'h00;
		ram[15'h12A] =  8'h00;
		ram[15'h12B] =  8'h00;
		ram[15'h12C] =  8'h00;
		ram[15'h12D] =  8'hFF;
		ram[15'h12E] =  8'hFF;
		ram[15'h12F] =  8'hFF;
		ram[15'h130] =  8'hFF;
		ram[15'h131] =  8'hFF;
		ram[15'h132] =  8'hFF;
		ram[15'h133] =  8'hD7;
		ram[15'h134] =  8'h00;
		ram[15'h135] =  8'hFF;
		ram[15'h136] =  8'hFF;
		ram[15'h137] =  8'hF8;
		ram[15'h138] =  8'hB4;
		ram[15'h139] =  8'hEA;
		ram[15'h13A] =  8'hA9;
		ram[15'h13B] =  8'h3C;
		ram[15'h13C] =  8'h61;
		ram[15'h13D] =  8'h64;
		ram[15'h13E] =  8'h63;
		ram[15'h13F] =  8'h2C;
		ram[15'h140] =  8'h73;
		ram[15'h141] =  8'h62;
		ram[15'h142] =  8'h63;
		ram[15'h143] =  8'h3E;
		ram[15'h144] =  8'h20;
		ram[15'h145] =  8'h68;
		ram[15'h146] =  8'h6C;
		ram[15'h147] =  8'h2C;
		ram[15'h148] =  8'h3C;
		ram[15'h149] =  8'h62;
		ram[15'h14A] =  8'h63;
		ram[15'h14B] =  8'h2C;
		ram[15'h14C] =  8'h64;
		ram[15'h14D] =  8'h65;
		ram[15'h14E] =  8'h2C;
		ram[15'h14F] =  8'h68;
		ram[15'h150] =  8'h6C;
		ram[15'h151] =  8'h2C;
		ram[15'h152] =  8'h73;
		ram[15'h153] =  8'h70;
		ram[15'h154] =  8'h3E;
		ram[15'h155] =  8'h2E;
		ram[15'h156] =  8'h2E;
		ram[15'h157] =  8'h2E;
		ram[15'h158] =  8'h2E;
		ram[15'h159] =  8'h24;
		ram[15'h15A] =  8'hC7;
		ram[15'h15B] =  8'h09;
		ram[15'h15C] =  8'h00;
		ram[15'h15D] =  8'h00;
		ram[15'h15E] =  8'h00;
		ram[15'h15F] =  8'hA5;
		ram[15'h160] =  8'hC4;
		ram[15'h161] =  8'hC7;
		ram[15'h162] =  8'hC4;
		ram[15'h163] =  8'h26;
		ram[15'h164] =  8'hD2;
		ram[15'h165] =  8'h50;
		ram[15'h166] =  8'hA0;
		ram[15'h167] =  8'hEA;
		ram[15'h168] =  8'h58;
		ram[15'h169] =  8'h66;
		ram[15'h16A] =  8'h85;
		ram[15'h16B] =  8'hC6;
		ram[15'h16C] =  8'hDE;
		ram[15'h16D] =  8'hC9;
		ram[15'h16E] =  8'h9B;
		ram[15'h16F] =  8'h30;
		ram[15'h170] =  8'h00;
		ram[15'h171] =  8'h00;
		ram[15'h172] =  8'h00;
		ram[15'h173] =  8'h00;
		ram[15'h174] =  8'h00;
		ram[15'h175] =  8'h00;
		ram[15'h176] =  8'h00;
		ram[15'h177] =  8'h00;
		ram[15'h178] =  8'h00;
		ram[15'h179] =  8'h21;
		ram[15'h17A] =  8'hF8;
		ram[15'h17B] =  8'h00;
		ram[15'h17C] =  8'h00;
		ram[15'h17D] =  8'h00;
		ram[15'h17E] =  8'h00;
		ram[15'h17F] =  8'h00;
		ram[15'h180] =  8'h00;
		ram[15'h181] =  8'h00;
		ram[15'h182] =  8'h00;
		ram[15'h183] =  8'h00;
		ram[15'h184] =  8'h00;
		ram[15'h185] =  8'h00;
		ram[15'h186] =  8'h00;
		ram[15'h187] =  8'h00;
		ram[15'h188] =  8'h00;
		ram[15'h189] =  8'h00;
		ram[15'h18A] =  8'h00;
		ram[15'h18B] =  8'h00;
		ram[15'h18C] =  8'h00;
		ram[15'h18D] =  8'hFF;
		ram[15'h18E] =  8'hFF;
		ram[15'h18F] =  8'hFF;
		ram[15'h190] =  8'hFF;
		ram[15'h191] =  8'hFF;
		ram[15'h192] =  8'hFF;
		ram[15'h193] =  8'hD7;
		ram[15'h194] =  8'h00;
		ram[15'h195] =  8'hFF;
		ram[15'h196] =  8'hFF;
		ram[15'h197] =  8'h89;
		ram[15'h198] =  8'hFD;
		ram[15'h199] =  8'hB6;
		ram[15'h19A] =  8'h35;
		ram[15'h19B] =  8'h61;
		ram[15'h19C] =  8'h64;
		ram[15'h19D] =  8'h64;
		ram[15'h19E] =  8'h20;
		ram[15'h19F] =  8'h68;
		ram[15'h1A0] =  8'h6C;
		ram[15'h1A1] =  8'h2C;
		ram[15'h1A2] =  8'h3C;
		ram[15'h1A3] =  8'h62;
		ram[15'h1A4] =  8'h63;
		ram[15'h1A5] =  8'h2C;
		ram[15'h1A6] =  8'h64;
		ram[15'h1A7] =  8'h65;
		ram[15'h1A8] =  8'h2C;
		ram[15'h1A9] =  8'h68;
		ram[15'h1AA] =  8'h6C;
		ram[15'h1AB] =  8'h2C;
		ram[15'h1AC] =  8'h73;
		ram[15'h1AD] =  8'h70;
		ram[15'h1AE] =  8'h3E;
		ram[15'h1AF] =  8'h2E;
		ram[15'h1B0] =  8'h2E;
		ram[15'h1B1] =  8'h2E;
		ram[15'h1B2] =  8'h2E;
		ram[15'h1B3] =  8'h2E;
		ram[15'h1B4] =  8'h2E;
		ram[15'h1B5] =  8'h2E;
		ram[15'h1B6] =  8'h2E;
		ram[15'h1B7] =  8'h2E;
		ram[15'h1B8] =  8'h2E;
		ram[15'h1B9] =  8'h24;
		ram[15'h1BA] =  8'hC7;
		ram[15'h1BB] =  8'hDD;
		ram[15'h1BC] =  8'h09;
		ram[15'h1BD] =  8'h00;
		ram[15'h1BE] =  8'h00;
		ram[15'h1BF] =  8'hAC;
		ram[15'h1C0] =  8'hDD;
		ram[15'h1C1] =  8'h94;
		ram[15'h1C2] =  8'hC2;
		ram[15'h1C3] =  8'h5B;
		ram[15'h1C4] =  8'h63;
		ram[15'h1C5] =  8'hD3;
		ram[15'h1C6] =  8'h33;
		ram[15'h1C7] =  8'h76;
		ram[15'h1C8] =  8'h6A;
		ram[15'h1C9] =  8'h20;
		ram[15'h1CA] =  8'hFA;
		ram[15'h1CB] =  8'h94;
		ram[15'h1CC] =  8'h68;
		ram[15'h1CD] =  8'hF5;
		ram[15'h1CE] =  8'h36;
		ram[15'h1CF] =  8'h00;
		ram[15'h1D0] =  8'h30;
		ram[15'h1D1] =  8'h00;
		ram[15'h1D2] =  8'h00;
		ram[15'h1D3] =  8'h00;
		ram[15'h1D4] =  8'h00;
		ram[15'h1D5] =  8'h00;
		ram[15'h1D6] =  8'h00;
		ram[15'h1D7] =  8'h21;
		ram[15'h1D8] =  8'hF8;
		ram[15'h1D9] =  8'h00;
		ram[15'h1DA] =  8'h00;
		ram[15'h1DB] =  8'h00;
		ram[15'h1DC] =  8'h00;
		ram[15'h1DD] =  8'h00;
		ram[15'h1DE] =  8'h00;
		ram[15'h1DF] =  8'h00;
		ram[15'h1E0] =  8'h00;
		ram[15'h1E1] =  8'h00;
		ram[15'h1E2] =  8'h00;
		ram[15'h1E3] =  8'h00;
		ram[15'h1E4] =  8'h00;
		ram[15'h1E5] =  8'h00;
		ram[15'h1E6] =  8'h00;
		ram[15'h1E7] =  8'h00;
		ram[15'h1E8] =  8'h00;
		ram[15'h1E9] =  8'h00;
		ram[15'h1EA] =  8'h00;
		ram[15'h1EB] =  8'hFF;
		ram[15'h1EC] =  8'hFF;
		ram[15'h1ED] =  8'h00;
		ram[15'h1EE] =  8'h00;
		ram[15'h1EF] =  8'hFF;
		ram[15'h1F0] =  8'hFF;
		ram[15'h1F1] =  8'hFF;
		ram[15'h1F2] =  8'hFF;
		ram[15'h1F3] =  8'hD7;
		ram[15'h1F4] =  8'h00;
		ram[15'h1F5] =  8'hFF;
		ram[15'h1F6] =  8'hFF;
		ram[15'h1F7] =  8'hC1;
		ram[15'h1F8] =  8'h33;
		ram[15'h1F9] =  8'h79;
		ram[15'h1FA] =  8'h0B;
		ram[15'h1FB] =  8'h61;
		ram[15'h1FC] =  8'h64;
		ram[15'h1FD] =  8'h64;
		ram[15'h1FE] =  8'h20;
		ram[15'h1FF] =  8'h69;
		ram[15'h200] =  8'h78;
		ram[15'h201] =  8'h2C;
		ram[15'h202] =  8'h3C;
		ram[15'h203] =  8'h62;
		ram[15'h204] =  8'h63;
		ram[15'h205] =  8'h2C;
		ram[15'h206] =  8'h64;
		ram[15'h207] =  8'h65;
		ram[15'h208] =  8'h2C;
		ram[15'h209] =  8'h69;
		ram[15'h20A] =  8'h78;
		ram[15'h20B] =  8'h2C;
		ram[15'h20C] =  8'h73;
		ram[15'h20D] =  8'h70;
		ram[15'h20E] =  8'h3E;
		ram[15'h20F] =  8'h2E;
		ram[15'h210] =  8'h2E;
		ram[15'h211] =  8'h2E;
		ram[15'h212] =  8'h2E;
		ram[15'h213] =  8'h2E;
		ram[15'h214] =  8'h2E;
		ram[15'h215] =  8'h2E;
		ram[15'h216] =  8'h2E;
		ram[15'h217] =  8'h2E;
		ram[15'h218] =  8'h2E;
		ram[15'h219] =  8'h24;
		ram[15'h21A] =  8'hC7;
		ram[15'h21B] =  8'hFD;
		ram[15'h21C] =  8'h09;
		ram[15'h21D] =  8'h00;
		ram[15'h21E] =  8'h00;
		ram[15'h21F] =  8'hC2;
		ram[15'h220] =  8'hC7;
		ram[15'h221] =  8'h07;
		ram[15'h222] =  8'hF4;
		ram[15'h223] =  8'hC1;
		ram[15'h224] =  8'h51;
		ram[15'h225] =  8'h96;
		ram[15'h226] =  8'h3E;
		ram[15'h227] =  8'hF4;
		ram[15'h228] =  8'h0B;
		ram[15'h229] =  8'h0F;
		ram[15'h22A] =  8'h51;
		ram[15'h22B] =  8'h92;
		ram[15'h22C] =  8'h1E;
		ram[15'h22D] =  8'hEA;
		ram[15'h22E] =  8'h71;
		ram[15'h22F] =  8'h00;
		ram[15'h230] =  8'h30;
		ram[15'h231] =  8'h00;
		ram[15'h232] =  8'h00;
		ram[15'h233] =  8'h00;
		ram[15'h234] =  8'h00;
		ram[15'h235] =  8'h21;
		ram[15'h236] =  8'hF8;
		ram[15'h237] =  8'h00;
		ram[15'h238] =  8'h00;
		ram[15'h239] =  8'h00;
		ram[15'h23A] =  8'h00;
		ram[15'h23B] =  8'h00;
		ram[15'h23C] =  8'h00;
		ram[15'h23D] =  8'h00;
		ram[15'h23E] =  8'h00;
		ram[15'h23F] =  8'h00;
		ram[15'h240] =  8'h00;
		ram[15'h241] =  8'h00;
		ram[15'h242] =  8'h00;
		ram[15'h243] =  8'h00;
		ram[15'h244] =  8'h00;
		ram[15'h245] =  8'h00;
		ram[15'h246] =  8'h00;
		ram[15'h247] =  8'h00;
		ram[15'h248] =  8'h00;
		ram[15'h249] =  8'hFF;
		ram[15'h24A] =  8'hFF;
		ram[15'h24B] =  8'h00;
		ram[15'h24C] =  8'h00;
		ram[15'h24D] =  8'h00;
		ram[15'h24E] =  8'h00;
		ram[15'h24F] =  8'hFF;
		ram[15'h250] =  8'hFF;
		ram[15'h251] =  8'hFF;
		ram[15'h252] =  8'hFF;
		ram[15'h253] =  8'hD7;
		ram[15'h254] =  8'h00;
		ram[15'h255] =  8'hFF;
		ram[15'h256] =  8'hFF;
		ram[15'h257] =  8'hE8;
		ram[15'h258] =  8'h81;
		ram[15'h259] =  8'h7B;
		ram[15'h25A] =  8'h9E;
		ram[15'h25B] =  8'h61;
		ram[15'h25C] =  8'h64;
		ram[15'h25D] =  8'h64;
		ram[15'h25E] =  8'h20;
		ram[15'h25F] =  8'h69;
		ram[15'h260] =  8'h79;
		ram[15'h261] =  8'h2C;
		ram[15'h262] =  8'h3C;
		ram[15'h263] =  8'h62;
		ram[15'h264] =  8'h63;
		ram[15'h265] =  8'h2C;
		ram[15'h266] =  8'h64;
		ram[15'h267] =  8'h65;
		ram[15'h268] =  8'h2C;
		ram[15'h269] =  8'h69;
		ram[15'h26A] =  8'h79;
		ram[15'h26B] =  8'h2C;
		ram[15'h26C] =  8'h73;
		ram[15'h26D] =  8'h70;
		ram[15'h26E] =  8'h3E;
		ram[15'h26F] =  8'h2E;
		ram[15'h270] =  8'h2E;
		ram[15'h271] =  8'h2E;
		ram[15'h272] =  8'h2E;
		ram[15'h273] =  8'h2E;
		ram[15'h274] =  8'h2E;
		ram[15'h275] =  8'h2E;
		ram[15'h276] =  8'h2E;
		ram[15'h277] =  8'h2E;
		ram[15'h278] =  8'h2E;
		ram[15'h279] =  8'h24;
		ram[15'h27A] =  8'hD7;
		ram[15'h27B] =  8'hC6;
		ram[15'h27C] =  8'h00;
		ram[15'h27D] =  8'h00;
		ram[15'h27E] =  8'h00;
		ram[15'h27F] =  8'h40;
		ram[15'h280] =  8'h91;
		ram[15'h281] =  8'h3C;
		ram[15'h282] =  8'h7E;
		ram[15'h283] =  8'h67;
		ram[15'h284] =  8'h7A;
		ram[15'h285] =  8'h6D;
		ram[15'h286] =  8'hDF;
		ram[15'h287] =  8'h61;
		ram[15'h288] =  8'h5B;
		ram[15'h289] =  8'h29;
		ram[15'h28A] =  8'h0B;
		ram[15'h28B] =  8'h10;
		ram[15'h28C] =  8'h66;
		ram[15'h28D] =  8'hB2;
		ram[15'h28E] =  8'h85;
		ram[15'h28F] =  8'h38;
		ram[15'h290] =  8'h00;
		ram[15'h291] =  8'h00;
		ram[15'h292] =  8'h00;
		ram[15'h293] =  8'h00;
		ram[15'h294] =  8'h00;
		ram[15'h295] =  8'h00;
		ram[15'h296] =  8'h00;
		ram[15'h297] =  8'h00;
		ram[15'h298] =  8'h00;
		ram[15'h299] =  8'h00;
		ram[15'h29A] =  8'h00;
		ram[15'h29B] =  8'h00;
		ram[15'h29C] =  8'h00;
		ram[15'h29D] =  8'h00;
		ram[15'h29E] =  8'h00;
		ram[15'h29F] =  8'h00;
		ram[15'h2A0] =  8'hFF;
		ram[15'h2A1] =  8'h00;
		ram[15'h2A2] =  8'h00;
		ram[15'h2A3] =  8'h00;
		ram[15'h2A4] =  8'hFF;
		ram[15'h2A5] =  8'h00;
		ram[15'h2A6] =  8'h00;
		ram[15'h2A7] =  8'h00;
		ram[15'h2A8] =  8'h00;
		ram[15'h2A9] =  8'h00;
		ram[15'h2AA] =  8'h00;
		ram[15'h2AB] =  8'h00;
		ram[15'h2AC] =  8'h00;
		ram[15'h2AD] =  8'h00;
		ram[15'h2AE] =  8'h00;
		ram[15'h2AF] =  8'h00;
		ram[15'h2B0] =  8'h00;
		ram[15'h2B1] =  8'h00;
		ram[15'h2B2] =  8'h00;
		ram[15'h2B3] =  8'hD7;
		ram[15'h2B4] =  8'h00;
		ram[15'h2B5] =  8'h00;
		ram[15'h2B6] =  8'h00;
		ram[15'h2B7] =  8'h48;
		ram[15'h2B8] =  8'h79;
		ram[15'h2B9] =  8'h93;
		ram[15'h2BA] =  8'h60;
		ram[15'h2BB] =  8'h61;
		ram[15'h2BC] =  8'h6C;
		ram[15'h2BD] =  8'h75;
		ram[15'h2BE] =  8'h6F;
		ram[15'h2BF] =  8'h70;
		ram[15'h2C0] =  8'h20;
		ram[15'h2C1] =  8'h61;
		ram[15'h2C2] =  8'h2C;
		ram[15'h2C3] =  8'h6E;
		ram[15'h2C4] =  8'h6E;
		ram[15'h2C5] =  8'h2E;
		ram[15'h2C6] =  8'h2E;
		ram[15'h2C7] =  8'h2E;
		ram[15'h2C8] =  8'h2E;
		ram[15'h2C9] =  8'h2E;
		ram[15'h2CA] =  8'h2E;
		ram[15'h2CB] =  8'h2E;
		ram[15'h2CC] =  8'h2E;
		ram[15'h2CD] =  8'h2E;
		ram[15'h2CE] =  8'h2E;
		ram[15'h2CF] =  8'h2E;
		ram[15'h2D0] =  8'h2E;
		ram[15'h2D1] =  8'h2E;
		ram[15'h2D2] =  8'h2E;
		ram[15'h2D3] =  8'h2E;
		ram[15'h2D4] =  8'h2E;
		ram[15'h2D5] =  8'h2E;
		ram[15'h2D6] =  8'h2E;
		ram[15'h2D7] =  8'h2E;
		ram[15'h2D8] =  8'h2E;
		ram[15'h2D9] =  8'h24;
		ram[15'h2DA] =  8'hD7;
		ram[15'h2DB] =  8'h80;
		ram[15'h2DC] =  8'h00;
		ram[15'h2DD] =  8'h00;
		ram[15'h2DE] =  8'h00;
		ram[15'h2DF] =  8'h3E;
		ram[15'h2E0] =  8'hC5;
		ram[15'h2E1] =  8'h3A;
		ram[15'h2E2] =  8'h57;
		ram[15'h2E3] =  8'h4D;
		ram[15'h2E4] =  8'h4C;
		ram[15'h2E5] =  8'h3A;
		ram[15'h2E6] =  8'h00;
		ram[15'h2E7] =  8'h09;
		ram[15'h2E8] =  8'hE3;
		ram[15'h2E9] =  8'h66;
		ram[15'h2EA] =  8'hA6;
		ram[15'h2EB] =  8'hD0;
		ram[15'h2EC] =  8'h3B;
		ram[15'h2ED] =  8'hBB;
		ram[15'h2EE] =  8'hAD;
		ram[15'h2EF] =  8'h3F;
		ram[15'h2F0] =  8'h00;
		ram[15'h2F1] =  8'h00;
		ram[15'h2F2] =  8'h00;
		ram[15'h2F3] =  8'h00;
		ram[15'h2F4] =  8'h00;
		ram[15'h2F5] =  8'h00;
		ram[15'h2F6] =  8'h00;
		ram[15'h2F7] =  8'h00;
		ram[15'h2F8] =  8'h00;
		ram[15'h2F9] =  8'h00;
		ram[15'h2FA] =  8'h00;
		ram[15'h2FB] =  8'h00;
		ram[15'h2FC] =  8'h00;
		ram[15'h2FD] =  8'h00;
		ram[15'h2FE] =  8'h00;
		ram[15'h2FF] =  8'h00;
		ram[15'h300] =  8'hFF;
		ram[15'h301] =  8'h00;
		ram[15'h302] =  8'h00;
		ram[15'h303] =  8'h00;
		ram[15'h304] =  8'h00;
		ram[15'h305] =  8'h00;
		ram[15'h306] =  8'h00;
		ram[15'h307] =  8'hFF;
		ram[15'h308] =  8'h00;
		ram[15'h309] =  8'h00;
		ram[15'h30A] =  8'h00;
		ram[15'h30B] =  8'h00;
		ram[15'h30C] =  8'h00;
		ram[15'h30D] =  8'h00;
		ram[15'h30E] =  8'h00;
		ram[15'h30F] =  8'hFF;
		ram[15'h310] =  8'hFF;
		ram[15'h311] =  8'hFF;
		ram[15'h312] =  8'hFF;
		ram[15'h313] =  8'hD7;
		ram[15'h314] =  8'h00;
		ram[15'h315] =  8'h00;
		ram[15'h316] =  8'h00;
		ram[15'h317] =  8'hFE;
		ram[15'h318] =  8'h43;
		ram[15'h319] =  8'hB0;
		ram[15'h31A] =  8'h16;
		ram[15'h31B] =  8'h61;
		ram[15'h31C] =  8'h6C;
		ram[15'h31D] =  8'h75;
		ram[15'h31E] =  8'h6F;
		ram[15'h31F] =  8'h70;
		ram[15'h320] =  8'h20;
		ram[15'h321] =  8'h61;
		ram[15'h322] =  8'h2C;
		ram[15'h323] =  8'h3C;
		ram[15'h324] =  8'h62;
		ram[15'h325] =  8'h2C;
		ram[15'h326] =  8'h63;
		ram[15'h327] =  8'h2C;
		ram[15'h328] =  8'h64;
		ram[15'h329] =  8'h2C;
		ram[15'h32A] =  8'h65;
		ram[15'h32B] =  8'h2C;
		ram[15'h32C] =  8'h68;
		ram[15'h32D] =  8'h2C;
		ram[15'h32E] =  8'h6C;
		ram[15'h32F] =  8'h2C;
		ram[15'h330] =  8'h28;
		ram[15'h331] =  8'h68;
		ram[15'h332] =  8'h6C;
		ram[15'h333] =  8'h29;
		ram[15'h334] =  8'h2C;
		ram[15'h335] =  8'h61;
		ram[15'h336] =  8'h3E;
		ram[15'h337] =  8'h2E;
		ram[15'h338] =  8'h2E;
		ram[15'h339] =  8'h24;
		ram[15'h33A] =  8'hD7;
		ram[15'h33B] =  8'hDD;
		ram[15'h33C] =  8'h84;
		ram[15'h33D] =  8'h00;
		ram[15'h33E] =  8'h00;
		ram[15'h33F] =  8'hF7;
		ram[15'h340] =  8'hD6;
		ram[15'h341] =  8'h6E;
		ram[15'h342] =  8'hC7;
		ram[15'h343] =  8'hCF;
		ram[15'h344] =  8'hAC;
		ram[15'h345] =  8'h47;
		ram[15'h346] =  8'h28;
		ram[15'h347] =  8'hDD;
		ram[15'h348] =  8'h22;
		ram[15'h349] =  8'h35;
		ram[15'h34A] =  8'hC0;
		ram[15'h34B] =  8'hC5;
		ram[15'h34C] =  8'h38;
		ram[15'h34D] =  8'h4B;
		ram[15'h34E] =  8'h23;
		ram[15'h34F] =  8'h20;
		ram[15'h350] =  8'h39;
		ram[15'h351] =  8'h00;
		ram[15'h352] =  8'h00;
		ram[15'h353] =  8'h00;
		ram[15'h354] =  8'h00;
		ram[15'h355] =  8'h00;
		ram[15'h356] =  8'h00;
		ram[15'h357] =  8'h00;
		ram[15'h358] =  8'h00;
		ram[15'h359] =  8'h00;
		ram[15'h35A] =  8'h00;
		ram[15'h35B] =  8'h00;
		ram[15'h35C] =  8'h00;
		ram[15'h35D] =  8'h00;
		ram[15'h35E] =  8'h00;
		ram[15'h35F] =  8'h00;
		ram[15'h360] =  8'hFF;
		ram[15'h361] =  8'h00;
		ram[15'h362] =  8'h00;
		ram[15'h363] =  8'h00;
		ram[15'h364] =  8'h00;
		ram[15'h365] =  8'h00;
		ram[15'h366] =  8'h00;
		ram[15'h367] =  8'hFF;
		ram[15'h368] =  8'h00;
		ram[15'h369] =  8'h00;
		ram[15'h36A] =  8'h00;
		ram[15'h36B] =  8'h00;
		ram[15'h36C] =  8'h00;
		ram[15'h36D] =  8'h00;
		ram[15'h36E] =  8'h00;
		ram[15'h36F] =  8'hFF;
		ram[15'h370] =  8'hFF;
		ram[15'h371] =  8'hFF;
		ram[15'h372] =  8'hFF;
		ram[15'h373] =  8'hD7;
		ram[15'h374] =  8'h00;
		ram[15'h375] =  8'h00;
		ram[15'h376] =  8'h00;
		ram[15'h377] =  8'hA4;
		ram[15'h378] =  8'h02;
		ram[15'h379] =  8'h6D;
		ram[15'h37A] =  8'h5A;
		ram[15'h37B] =  8'h61;
		ram[15'h37C] =  8'h6C;
		ram[15'h37D] =  8'h75;
		ram[15'h37E] =  8'h6F;
		ram[15'h37F] =  8'h70;
		ram[15'h380] =  8'h20;
		ram[15'h381] =  8'h61;
		ram[15'h382] =  8'h2C;
		ram[15'h383] =  8'h3C;
		ram[15'h384] =  8'h69;
		ram[15'h385] =  8'h78;
		ram[15'h386] =  8'h68;
		ram[15'h387] =  8'h2C;
		ram[15'h388] =  8'h69;
		ram[15'h389] =  8'h78;
		ram[15'h38A] =  8'h6C;
		ram[15'h38B] =  8'h2C;
		ram[15'h38C] =  8'h69;
		ram[15'h38D] =  8'h79;
		ram[15'h38E] =  8'h68;
		ram[15'h38F] =  8'h2C;
		ram[15'h390] =  8'h69;
		ram[15'h391] =  8'h79;
		ram[15'h392] =  8'h6C;
		ram[15'h393] =  8'h3E;
		ram[15'h394] =  8'h2E;
		ram[15'h395] =  8'h2E;
		ram[15'h396] =  8'h2E;
		ram[15'h397] =  8'h2E;
		ram[15'h398] =  8'h2E;
		ram[15'h399] =  8'h24;
		ram[15'h39A] =  8'hD7;
		ram[15'h39B] =  8'hDD;
		ram[15'h39C] =  8'h86;
		ram[15'h39D] =  8'h01;
		ram[15'h39E] =  8'h00;
		ram[15'h39F] =  8'hB7;
		ram[15'h3A0] =  8'h90;
		ram[15'h3A1] =  8'h39;
		ram[15'h3A2] =  8'h00;
		ram[15'h3A3] =  8'h39;
		ram[15'h3A4] =  8'h00;
		ram[15'h3A5] =  8'hFD;
		ram[15'h3A6] =  8'h32;
		ram[15'h3A7] =  8'h6E;
		ram[15'h3A8] =  8'h40;
		ram[15'h3A9] =  8'hDC;
		ram[15'h3AA] =  8'hC1;
		ram[15'h3AB] =  8'h45;
		ram[15'h3AC] =  8'h6E;
		ram[15'h3AD] =  8'hFA;
		ram[15'h3AE] =  8'hE5;
		ram[15'h3AF] =  8'h20;
		ram[15'h3B0] =  8'h38;
		ram[15'h3B1] =  8'h00;
		ram[15'h3B2] =  8'h00;
		ram[15'h3B3] =  8'h00;
		ram[15'h3B4] =  8'h00;
		ram[15'h3B5] =  8'h01;
		ram[15'h3B6] =  8'h00;
		ram[15'h3B7] =  8'h01;
		ram[15'h3B8] =  8'h00;
		ram[15'h3B9] =  8'h00;
		ram[15'h3BA] =  8'h00;
		ram[15'h3BB] =  8'h00;
		ram[15'h3BC] =  8'h00;
		ram[15'h3BD] =  8'h00;
		ram[15'h3BE] =  8'h00;
		ram[15'h3BF] =  8'h00;
		ram[15'h3C0] =  8'hFF;
		ram[15'h3C1] =  8'h00;
		ram[15'h3C2] =  8'h00;
		ram[15'h3C3] =  8'h00;
		ram[15'h3C4] =  8'h00;
		ram[15'h3C5] =  8'h00;
		ram[15'h3C6] =  8'h00;
		ram[15'h3C7] =  8'hFF;
		ram[15'h3C8] =  8'h00;
		ram[15'h3C9] =  8'h00;
		ram[15'h3CA] =  8'h00;
		ram[15'h3CB] =  8'h00;
		ram[15'h3CC] =  8'h00;
		ram[15'h3CD] =  8'h00;
		ram[15'h3CE] =  8'h00;
		ram[15'h3CF] =  8'h00;
		ram[15'h3D0] =  8'h00;
		ram[15'h3D1] =  8'h00;
		ram[15'h3D2] =  8'h00;
		ram[15'h3D3] =  8'hD7;
		ram[15'h3D4] =  8'h00;
		ram[15'h3D5] =  8'h00;
		ram[15'h3D6] =  8'h00;
		ram[15'h3D7] =  8'hE8;
		ram[15'h3D8] =  8'h49;
		ram[15'h3D9] =  8'h67;
		ram[15'h3DA] =  8'h6E;
		ram[15'h3DB] =  8'h61;
		ram[15'h3DC] =  8'h6C;
		ram[15'h3DD] =  8'h75;
		ram[15'h3DE] =  8'h6F;
		ram[15'h3DF] =  8'h70;
		ram[15'h3E0] =  8'h20;
		ram[15'h3E1] =  8'h61;
		ram[15'h3E2] =  8'h2C;
		ram[15'h3E3] =  8'h28;
		ram[15'h3E4] =  8'h3C;
		ram[15'h3E5] =  8'h69;
		ram[15'h3E6] =  8'h78;
		ram[15'h3E7] =  8'h2C;
		ram[15'h3E8] =  8'h69;
		ram[15'h3E9] =  8'h79;
		ram[15'h3EA] =  8'h3E;
		ram[15'h3EB] =  8'h2B;
		ram[15'h3EC] =  8'h31;
		ram[15'h3ED] =  8'h29;
		ram[15'h3EE] =  8'h2E;
		ram[15'h3EF] =  8'h2E;
		ram[15'h3F0] =  8'h2E;
		ram[15'h3F1] =  8'h2E;
		ram[15'h3F2] =  8'h2E;
		ram[15'h3F3] =  8'h2E;
		ram[15'h3F4] =  8'h2E;
		ram[15'h3F5] =  8'h2E;
		ram[15'h3F6] =  8'h2E;
		ram[15'h3F7] =  8'h2E;
		ram[15'h3F8] =  8'h2E;
		ram[15'h3F9] =  8'h24;
		ram[15'h3FA] =  8'h53;
		ram[15'h3FB] =  8'hDD;
		ram[15'h3FC] =  8'hCB;
		ram[15'h3FD] =  8'h01;
		ram[15'h3FE] =  8'h46;
		ram[15'h3FF] =  8'h75;
		ram[15'h400] =  8'h20;
		ram[15'h401] =  8'h39;
		ram[15'h402] =  8'h00;
		ram[15'h403] =  8'h39;
		ram[15'h404] =  8'h00;
		ram[15'h405] =  8'hFC;
		ram[15'h406] =  8'h3C;
		ram[15'h407] =  8'h9A;
		ram[15'h408] =  8'hA7;
		ram[15'h409] =  8'h74;
		ram[15'h40A] =  8'h3D;
		ram[15'h40B] =  8'h51;
		ram[15'h40C] =  8'h27;
		ram[15'h40D] =  8'h14;
		ram[15'h40E] =  8'hCA;
		ram[15'h40F] =  8'h20;
		ram[15'h410] =  8'h00;
		ram[15'h411] =  8'h00;
		ram[15'h412] =  8'h38;
		ram[15'h413] =  8'h00;
		ram[15'h414] =  8'h00;
		ram[15'h415] =  8'h00;
		ram[15'h416] =  8'h00;
		ram[15'h417] =  8'h00;
		ram[15'h418] =  8'h00;
		ram[15'h419] =  8'h00;
		ram[15'h41A] =  8'h00;
		ram[15'h41B] =  8'h00;
		ram[15'h41C] =  8'h00;
		ram[15'h41D] =  8'h00;
		ram[15'h41E] =  8'h00;
		ram[15'h41F] =  8'h53;
		ram[15'h420] =  8'h00;
		ram[15'h421] =  8'h00;
		ram[15'h422] =  8'h00;
		ram[15'h423] =  8'h00;
		ram[15'h424] =  8'h00;
		ram[15'h425] =  8'h00;
		ram[15'h426] =  8'h00;
		ram[15'h427] =  8'hFF;
		ram[15'h428] =  8'h00;
		ram[15'h429] =  8'h00;
		ram[15'h42A] =  8'h00;
		ram[15'h42B] =  8'h00;
		ram[15'h42C] =  8'h00;
		ram[15'h42D] =  8'h00;
		ram[15'h42E] =  8'h00;
		ram[15'h42F] =  8'h00;
		ram[15'h430] =  8'h00;
		ram[15'h431] =  8'h00;
		ram[15'h432] =  8'h00;
		ram[15'h433] =  8'h00;
		ram[15'h434] =  8'h00;
		ram[15'h435] =  8'h00;
		ram[15'h436] =  8'h00;
		ram[15'h437] =  8'hA8;
		ram[15'h438] =  8'hEE;
		ram[15'h439] =  8'h08;
		ram[15'h43A] =  8'h67;
		ram[15'h43B] =  8'h62;
		ram[15'h43C] =  8'h69;
		ram[15'h43D] =  8'h74;
		ram[15'h43E] =  8'h20;
		ram[15'h43F] =  8'h6E;
		ram[15'h440] =  8'h2C;
		ram[15'h441] =  8'h28;
		ram[15'h442] =  8'h3C;
		ram[15'h443] =  8'h69;
		ram[15'h444] =  8'h78;
		ram[15'h445] =  8'h2C;
		ram[15'h446] =  8'h69;
		ram[15'h447] =  8'h79;
		ram[15'h448] =  8'h3E;
		ram[15'h449] =  8'h2B;
		ram[15'h44A] =  8'h31;
		ram[15'h44B] =  8'h29;
		ram[15'h44C] =  8'h2E;
		ram[15'h44D] =  8'h2E;
		ram[15'h44E] =  8'h2E;
		ram[15'h44F] =  8'h2E;
		ram[15'h450] =  8'h2E;
		ram[15'h451] =  8'h2E;
		ram[15'h452] =  8'h2E;
		ram[15'h453] =  8'h2E;
		ram[15'h454] =  8'h2E;
		ram[15'h455] =  8'h2E;
		ram[15'h456] =  8'h2E;
		ram[15'h457] =  8'h2E;
		ram[15'h458] =  8'h2E;
		ram[15'h459] =  8'h24;
		ram[15'h45A] =  8'h53;
		ram[15'h45B] =  8'hCB;
		ram[15'h45C] =  8'h40;
		ram[15'h45D] =  8'h00;
		ram[15'h45E] =  8'h00;
		ram[15'h45F] =  8'hF1;
		ram[15'h460] =  8'h3E;
		ram[15'h461] =  8'hFC;
		ram[15'h462] =  8'h9D;
		ram[15'h463] =  8'hCC;
		ram[15'h464] =  8'h7A;
		ram[15'h465] =  8'h3A;
		ram[15'h466] =  8'h00;
		ram[15'h467] =  8'h61;
		ram[15'h468] =  8'hBE;
		ram[15'h469] =  8'h86;
		ram[15'h46A] =  8'h7A;
		ram[15'h46B] =  8'h50;
		ram[15'h46C] =  8'h24;
		ram[15'h46D] =  8'h98;
		ram[15'h46E] =  8'h19;
		ram[15'h46F] =  8'h00;
		ram[15'h470] =  8'h3F;
		ram[15'h471] =  8'h00;
		ram[15'h472] =  8'h00;
		ram[15'h473] =  8'h00;
		ram[15'h474] =  8'h00;
		ram[15'h475] =  8'h00;
		ram[15'h476] =  8'h00;
		ram[15'h477] =  8'h00;
		ram[15'h478] =  8'h00;
		ram[15'h479] =  8'h00;
		ram[15'h47A] =  8'h00;
		ram[15'h47B] =  8'h00;
		ram[15'h47C] =  8'h00;
		ram[15'h47D] =  8'h00;
		ram[15'h47E] =  8'h00;
		ram[15'h47F] =  8'h53;
		ram[15'h480] =  8'h00;
		ram[15'h481] =  8'h00;
		ram[15'h482] =  8'h00;
		ram[15'h483] =  8'h00;
		ram[15'h484] =  8'h00;
		ram[15'h485] =  8'h00;
		ram[15'h486] =  8'h00;
		ram[15'h487] =  8'hFF;
		ram[15'h488] =  8'h00;
		ram[15'h489] =  8'h00;
		ram[15'h48A] =  8'h00;
		ram[15'h48B] =  8'h00;
		ram[15'h48C] =  8'h00;
		ram[15'h48D] =  8'h00;
		ram[15'h48E] =  8'h00;
		ram[15'h48F] =  8'hFF;
		ram[15'h490] =  8'hFF;
		ram[15'h491] =  8'hFF;
		ram[15'h492] =  8'hFF;
		ram[15'h493] =  8'h00;
		ram[15'h494] =  8'hFF;
		ram[15'h495] =  8'h00;
		ram[15'h496] =  8'h00;
		ram[15'h497] =  8'h7B;
		ram[15'h498] =  8'h55;
		ram[15'h499] =  8'hE6;
		ram[15'h49A] =  8'hC8;
		ram[15'h49B] =  8'h62;
		ram[15'h49C] =  8'h69;
		ram[15'h49D] =  8'h74;
		ram[15'h49E] =  8'h20;
		ram[15'h49F] =  8'h6E;
		ram[15'h4A0] =  8'h2C;
		ram[15'h4A1] =  8'h3C;
		ram[15'h4A2] =  8'h62;
		ram[15'h4A3] =  8'h2C;
		ram[15'h4A4] =  8'h63;
		ram[15'h4A5] =  8'h2C;
		ram[15'h4A6] =  8'h64;
		ram[15'h4A7] =  8'h2C;
		ram[15'h4A8] =  8'h65;
		ram[15'h4A9] =  8'h2C;
		ram[15'h4AA] =  8'h68;
		ram[15'h4AB] =  8'h2C;
		ram[15'h4AC] =  8'h6C;
		ram[15'h4AD] =  8'h2C;
		ram[15'h4AE] =  8'h28;
		ram[15'h4AF] =  8'h68;
		ram[15'h4B0] =  8'h6C;
		ram[15'h4B1] =  8'h29;
		ram[15'h4B2] =  8'h2C;
		ram[15'h4B3] =  8'h61;
		ram[15'h4B4] =  8'h3E;
		ram[15'h4B5] =  8'h2E;
		ram[15'h4B6] =  8'h2E;
		ram[15'h4B7] =  8'h2E;
		ram[15'h4B8] =  8'h2E;
		ram[15'h4B9] =  8'h24;
		ram[15'h4BA] =  8'hD7;
		ram[15'h4BB] =  8'hED;
		ram[15'h4BC] =  8'hA9;
		ram[15'h4BD] =  8'h00;
		ram[15'h4BE] =  8'h00;
		ram[15'h4BF] =  8'hB6;
		ram[15'h4C0] =  8'hC7;
		ram[15'h4C1] =  8'hB4;
		ram[15'h4C2] =  8'h72;
		ram[15'h4C3] =  8'hF6;
		ram[15'h4C4] =  8'h18;
		ram[15'h4C5] =  8'h4B;
		ram[15'h4C6] =  8'h00;
		ram[15'h4C7] =  8'hBD;
		ram[15'h4C8] =  8'h8D;
		ram[15'h4C9] =  8'h01;
		ram[15'h4CA] =  8'h00;
		ram[15'h4CB] =  8'hC0;
		ram[15'h4CC] =  8'h30;
		ram[15'h4CD] =  8'hA3;
		ram[15'h4CE] =  8'h94;
		ram[15'h4CF] =  8'h00;
		ram[15'h4D0] =  8'h10;
		ram[15'h4D1] =  8'h00;
		ram[15'h4D2] =  8'h00;
		ram[15'h4D3] =  8'h00;
		ram[15'h4D4] =  8'h00;
		ram[15'h4D5] =  8'h00;
		ram[15'h4D6] =  8'h00;
		ram[15'h4D7] =  8'h00;
		ram[15'h4D8] =  8'h00;
		ram[15'h4D9] =  8'h00;
		ram[15'h4DA] =  8'h00;
		ram[15'h4DB] =  8'h00;
		ram[15'h4DC] =  8'h00;
		ram[15'h4DD] =  8'h0A;
		ram[15'h4DE] =  8'h00;
		ram[15'h4DF] =  8'h00;
		ram[15'h4E0] =  8'hFF;
		ram[15'h4E1] =  8'h00;
		ram[15'h4E2] =  8'h00;
		ram[15'h4E3] =  8'h00;
		ram[15'h4E4] =  8'h00;
		ram[15'h4E5] =  8'h00;
		ram[15'h4E6] =  8'h00;
		ram[15'h4E7] =  8'h00;
		ram[15'h4E8] =  8'h00;
		ram[15'h4E9] =  8'h00;
		ram[15'h4EA] =  8'h00;
		ram[15'h4EB] =  8'h00;
		ram[15'h4EC] =  8'h00;
		ram[15'h4ED] =  8'h00;
		ram[15'h4EE] =  8'h00;
		ram[15'h4EF] =  8'h00;
		ram[15'h4F0] =  8'h00;
		ram[15'h4F1] =  8'h00;
		ram[15'h4F2] =  8'h00;
		ram[15'h4F3] =  8'hD7;
		ram[15'h4F4] =  8'h00;
		ram[15'h4F5] =  8'h00;
		ram[15'h4F6] =  8'h00;
		ram[15'h4F7] =  8'hA8;
		ram[15'h4F8] =  8'h7E;
		ram[15'h4F9] =  8'h6C;
		ram[15'h4FA] =  8'hFA;
		ram[15'h4FB] =  8'h63;
		ram[15'h4FC] =  8'h70;
		ram[15'h4FD] =  8'h64;
		ram[15'h4FE] =  8'h3C;
		ram[15'h4FF] =  8'h72;
		ram[15'h500] =  8'h3E;
		ram[15'h501] =  8'h2E;
		ram[15'h502] =  8'h2E;
		ram[15'h503] =  8'h2E;
		ram[15'h504] =  8'h2E;
		ram[15'h505] =  8'h2E;
		ram[15'h506] =  8'h2E;
		ram[15'h507] =  8'h2E;
		ram[15'h508] =  8'h2E;
		ram[15'h509] =  8'h2E;
		ram[15'h50A] =  8'h2E;
		ram[15'h50B] =  8'h2E;
		ram[15'h50C] =  8'h2E;
		ram[15'h50D] =  8'h2E;
		ram[15'h50E] =  8'h2E;
		ram[15'h50F] =  8'h2E;
		ram[15'h510] =  8'h2E;
		ram[15'h511] =  8'h2E;
		ram[15'h512] =  8'h2E;
		ram[15'h513] =  8'h2E;
		ram[15'h514] =  8'h2E;
		ram[15'h515] =  8'h2E;
		ram[15'h516] =  8'h2E;
		ram[15'h517] =  8'h2E;
		ram[15'h518] =  8'h2E;
		ram[15'h519] =  8'h24;
		ram[15'h51A] =  8'hD7;
		ram[15'h51B] =  8'hED;
		ram[15'h51C] =  8'hA1;
		ram[15'h51D] =  8'h00;
		ram[15'h51E] =  8'h00;
		ram[15'h51F] =  8'h48;
		ram[15'h520] =  8'h4D;
		ram[15'h521] =  8'h4A;
		ram[15'h522] =  8'hAF;
		ram[15'h523] =  8'h6B;
		ram[15'h524] =  8'h90;
		ram[15'h525] =  8'h3A;
		ram[15'h526] =  8'h00;
		ram[15'h527] =  8'h71;
		ram[15'h528] =  8'h4E;
		ram[15'h529] =  8'h01;
		ram[15'h52A] =  8'h00;
		ram[15'h52B] =  8'h93;
		ram[15'h52C] =  8'h6A;
		ram[15'h52D] =  8'h7C;
		ram[15'h52E] =  8'h90;
		ram[15'h52F] =  8'h00;
		ram[15'h530] =  8'h10;
		ram[15'h531] =  8'h00;
		ram[15'h532] =  8'h00;
		ram[15'h533] =  8'h00;
		ram[15'h534] =  8'h00;
		ram[15'h535] =  8'h00;
		ram[15'h536] =  8'h00;
		ram[15'h537] =  8'h00;
		ram[15'h538] =  8'h00;
		ram[15'h539] =  8'h00;
		ram[15'h53A] =  8'h00;
		ram[15'h53B] =  8'h00;
		ram[15'h53C] =  8'h00;
		ram[15'h53D] =  8'h0A;
		ram[15'h53E] =  8'h00;
		ram[15'h53F] =  8'h00;
		ram[15'h540] =  8'hFF;
		ram[15'h541] =  8'h00;
		ram[15'h542] =  8'h00;
		ram[15'h543] =  8'h00;
		ram[15'h544] =  8'h00;
		ram[15'h545] =  8'h00;
		ram[15'h546] =  8'h00;
		ram[15'h547] =  8'h00;
		ram[15'h548] =  8'h00;
		ram[15'h549] =  8'h00;
		ram[15'h54A] =  8'h00;
		ram[15'h54B] =  8'h00;
		ram[15'h54C] =  8'h00;
		ram[15'h54D] =  8'h00;
		ram[15'h54E] =  8'h00;
		ram[15'h54F] =  8'h00;
		ram[15'h550] =  8'h00;
		ram[15'h551] =  8'h00;
		ram[15'h552] =  8'h00;
		ram[15'h553] =  8'hD7;
		ram[15'h554] =  8'h00;
		ram[15'h555] =  8'h00;
		ram[15'h556] =  8'h00;
		ram[15'h557] =  8'h06;
		ram[15'h558] =  8'hDE;
		ram[15'h559] =  8'hB3;
		ram[15'h55A] =  8'h56;
		ram[15'h55B] =  8'h63;
		ram[15'h55C] =  8'h70;
		ram[15'h55D] =  8'h69;
		ram[15'h55E] =  8'h3C;
		ram[15'h55F] =  8'h72;
		ram[15'h560] =  8'h3E;
		ram[15'h561] =  8'h2E;
		ram[15'h562] =  8'h2E;
		ram[15'h563] =  8'h2E;
		ram[15'h564] =  8'h2E;
		ram[15'h565] =  8'h2E;
		ram[15'h566] =  8'h2E;
		ram[15'h567] =  8'h2E;
		ram[15'h568] =  8'h2E;
		ram[15'h569] =  8'h2E;
		ram[15'h56A] =  8'h2E;
		ram[15'h56B] =  8'h2E;
		ram[15'h56C] =  8'h2E;
		ram[15'h56D] =  8'h2E;
		ram[15'h56E] =  8'h2E;
		ram[15'h56F] =  8'h2E;
		ram[15'h570] =  8'h2E;
		ram[15'h571] =  8'h2E;
		ram[15'h572] =  8'h2E;
		ram[15'h573] =  8'h2E;
		ram[15'h574] =  8'h2E;
		ram[15'h575] =  8'h2E;
		ram[15'h576] =  8'h2E;
		ram[15'h577] =  8'h2E;
		ram[15'h578] =  8'h2E;
		ram[15'h579] =  8'h24;
		ram[15'h57A] =  8'hD7;
		ram[15'h57B] =  8'h27;
		ram[15'h57C] =  8'h00;
		ram[15'h57D] =  8'h00;
		ram[15'h57E] =  8'h00;
		ram[15'h57F] =  8'h41;
		ram[15'h580] =  8'h21;
		ram[15'h581] =  8'hFA;
		ram[15'h582] =  8'h09;
		ram[15'h583] =  8'h60;
		ram[15'h584] =  8'h1D;
		ram[15'h585] =  8'h59;
		ram[15'h586] =  8'hA5;
		ram[15'h587] =  8'h5B;
		ram[15'h588] =  8'h8D;
		ram[15'h589] =  8'h79;
		ram[15'h58A] =  8'h90;
		ram[15'h58B] =  8'h04;
		ram[15'h58C] =  8'h8E;
		ram[15'h58D] =  8'h9D;
		ram[15'h58E] =  8'h29;
		ram[15'h58F] =  8'h18;
		ram[15'h590] =  8'h00;
		ram[15'h591] =  8'h00;
		ram[15'h592] =  8'h00;
		ram[15'h593] =  8'h00;
		ram[15'h594] =  8'h00;
		ram[15'h595] =  8'h00;
		ram[15'h596] =  8'h00;
		ram[15'h597] =  8'h00;
		ram[15'h598] =  8'h00;
		ram[15'h599] =  8'h00;
		ram[15'h59A] =  8'h00;
		ram[15'h59B] =  8'h00;
		ram[15'h59C] =  8'h00;
		ram[15'h59D] =  8'h00;
		ram[15'h59E] =  8'h00;
		ram[15'h59F] =  8'hD7;
		ram[15'h5A0] =  8'hFF;
		ram[15'h5A1] =  8'h00;
		ram[15'h5A2] =  8'h00;
		ram[15'h5A3] =  8'h00;
		ram[15'h5A4] =  8'h00;
		ram[15'h5A5] =  8'h00;
		ram[15'h5A6] =  8'h00;
		ram[15'h5A7] =  8'h00;
		ram[15'h5A8] =  8'h00;
		ram[15'h5A9] =  8'h00;
		ram[15'h5AA] =  8'h00;
		ram[15'h5AB] =  8'h00;
		ram[15'h5AC] =  8'h00;
		ram[15'h5AD] =  8'h00;
		ram[15'h5AE] =  8'h00;
		ram[15'h5AF] =  8'h00;
		ram[15'h5B0] =  8'h00;
		ram[15'h5B1] =  8'h00;
		ram[15'h5B2] =  8'h00;
		ram[15'h5B3] =  8'h00;
		ram[15'h5B4] =  8'h00;
		ram[15'h5B5] =  8'h00;
		ram[15'h5B6] =  8'h00;
		ram[15'h5B7] =  8'h9B;
		ram[15'h5B8] =  8'h4B;
		ram[15'h5B9] =  8'hA6;
		ram[15'h5BA] =  8'h75;
		ram[15'h5BB] =  8'h3C;
		ram[15'h5BC] =  8'h64;
		ram[15'h5BD] =  8'h61;
		ram[15'h5BE] =  8'h61;
		ram[15'h5BF] =  8'h2C;
		ram[15'h5C0] =  8'h63;
		ram[15'h5C1] =  8'h70;
		ram[15'h5C2] =  8'h6C;
		ram[15'h5C3] =  8'h2C;
		ram[15'h5C4] =  8'h73;
		ram[15'h5C5] =  8'h63;
		ram[15'h5C6] =  8'h66;
		ram[15'h5C7] =  8'h2C;
		ram[15'h5C8] =  8'h63;
		ram[15'h5C9] =  8'h63;
		ram[15'h5CA] =  8'h66;
		ram[15'h5CB] =  8'h3E;
		ram[15'h5CC] =  8'h2E;
		ram[15'h5CD] =  8'h2E;
		ram[15'h5CE] =  8'h2E;
		ram[15'h5CF] =  8'h2E;
		ram[15'h5D0] =  8'h2E;
		ram[15'h5D1] =  8'h2E;
		ram[15'h5D2] =  8'h2E;
		ram[15'h5D3] =  8'h2E;
		ram[15'h5D4] =  8'h2E;
		ram[15'h5D5] =  8'h2E;
		ram[15'h5D6] =  8'h2E;
		ram[15'h5D7] =  8'h2E;
		ram[15'h5D8] =  8'h2E;
		ram[15'h5D9] =  8'h24;
		ram[15'h5DA] =  8'hD7;
		ram[15'h5DB] =  8'h3C;
		ram[15'h5DC] =  8'h00;
		ram[15'h5DD] =  8'h00;
		ram[15'h5DE] =  8'h00;
		ram[15'h5DF] =  8'hDF;
		ram[15'h5E0] =  8'h4A;
		ram[15'h5E1] =  8'hD8;
		ram[15'h5E2] =  8'hD5;
		ram[15'h5E3] =  8'h98;
		ram[15'h5E4] =  8'hE5;
		ram[15'h5E5] =  8'h2B;
		ram[15'h5E6] =  8'h8A;
		ram[15'h5E7] =  8'hB0;
		ram[15'h5E8] =  8'hA7;
		ram[15'h5E9] =  8'h1B;
		ram[15'h5EA] =  8'h43;
		ram[15'h5EB] =  8'h44;
		ram[15'h5EC] =  8'h5A;
		ram[15'h5ED] =  8'h30;
		ram[15'h5EE] =  8'hD0;
		ram[15'h5EF] =  8'h01;
		ram[15'h5F0] =  8'h00;
		ram[15'h5F1] =  8'h00;
		ram[15'h5F2] =  8'h00;
		ram[15'h5F3] =  8'h00;
		ram[15'h5F4] =  8'h00;
		ram[15'h5F5] =  8'h00;
		ram[15'h5F6] =  8'h00;
		ram[15'h5F7] =  8'h00;
		ram[15'h5F8] =  8'h00;
		ram[15'h5F9] =  8'h00;
		ram[15'h5FA] =  8'h00;
		ram[15'h5FB] =  8'h00;
		ram[15'h5FC] =  8'h00;
		ram[15'h5FD] =  8'h00;
		ram[15'h5FE] =  8'h00;
		ram[15'h5FF] =  8'h00;
		ram[15'h600] =  8'hFF;
		ram[15'h601] =  8'h00;
		ram[15'h602] =  8'h00;
		ram[15'h603] =  8'h00;
		ram[15'h604] =  8'h00;
		ram[15'h605] =  8'h00;
		ram[15'h606] =  8'h00;
		ram[15'h607] =  8'h00;
		ram[15'h608] =  8'h00;
		ram[15'h609] =  8'h00;
		ram[15'h60A] =  8'h00;
		ram[15'h60B] =  8'h00;
		ram[15'h60C] =  8'h00;
		ram[15'h60D] =  8'h00;
		ram[15'h60E] =  8'h00;
		ram[15'h60F] =  8'h00;
		ram[15'h610] =  8'h00;
		ram[15'h611] =  8'h00;
		ram[15'h612] =  8'h00;
		ram[15'h613] =  8'hD7;
		ram[15'h614] =  8'h00;
		ram[15'h615] =  8'h00;
		ram[15'h616] =  8'h00;
		ram[15'h617] =  8'hD1;
		ram[15'h618] =  8'h88;
		ram[15'h619] =  8'h15;
		ram[15'h61A] =  8'hA4;
		ram[15'h61B] =  8'h3C;
		ram[15'h61C] =  8'h69;
		ram[15'h61D] =  8'h6E;
		ram[15'h61E] =  8'h63;
		ram[15'h61F] =  8'h2C;
		ram[15'h620] =  8'h64;
		ram[15'h621] =  8'h65;
		ram[15'h622] =  8'h63;
		ram[15'h623] =  8'h3E;
		ram[15'h624] =  8'h20;
		ram[15'h625] =  8'h61;
		ram[15'h626] =  8'h2E;
		ram[15'h627] =  8'h2E;
		ram[15'h628] =  8'h2E;
		ram[15'h629] =  8'h2E;
		ram[15'h62A] =  8'h2E;
		ram[15'h62B] =  8'h2E;
		ram[15'h62C] =  8'h2E;
		ram[15'h62D] =  8'h2E;
		ram[15'h62E] =  8'h2E;
		ram[15'h62F] =  8'h2E;
		ram[15'h630] =  8'h2E;
		ram[15'h631] =  8'h2E;
		ram[15'h632] =  8'h2E;
		ram[15'h633] =  8'h2E;
		ram[15'h634] =  8'h2E;
		ram[15'h635] =  8'h2E;
		ram[15'h636] =  8'h2E;
		ram[15'h637] =  8'h2E;
		ram[15'h638] =  8'h2E;
		ram[15'h639] =  8'h24;
		ram[15'h63A] =  8'hD7;
		ram[15'h63B] =  8'h04;
		ram[15'h63C] =  8'h00;
		ram[15'h63D] =  8'h00;
		ram[15'h63E] =  8'h00;
		ram[15'h63F] =  8'h23;
		ram[15'h640] =  8'hD6;
		ram[15'h641] =  8'h2D;
		ram[15'h642] =  8'h43;
		ram[15'h643] =  8'h61;
		ram[15'h644] =  8'h7A;
		ram[15'h645] =  8'h80;
		ram[15'h646] =  8'h81;
		ram[15'h647] =  8'h86;
		ram[15'h648] =  8'h5A;
		ram[15'h649] =  8'h85;
		ram[15'h64A] =  8'h1E;
		ram[15'h64B] =  8'h86;
		ram[15'h64C] =  8'h58;
		ram[15'h64D] =  8'hBB;
		ram[15'h64E] =  8'h9B;
		ram[15'h64F] =  8'h01;
		ram[15'h650] =  8'h00;
		ram[15'h651] =  8'h00;
		ram[15'h652] =  8'h00;
		ram[15'h653] =  8'h00;
		ram[15'h654] =  8'h00;
		ram[15'h655] =  8'h00;
		ram[15'h656] =  8'h00;
		ram[15'h657] =  8'h00;
		ram[15'h658] =  8'h00;
		ram[15'h659] =  8'h00;
		ram[15'h65A] =  8'h00;
		ram[15'h65B] =  8'h00;
		ram[15'h65C] =  8'h00;
		ram[15'h65D] =  8'h00;
		ram[15'h65E] =  8'hFF;
		ram[15'h65F] =  8'h00;
		ram[15'h660] =  8'h00;
		ram[15'h661] =  8'h00;
		ram[15'h662] =  8'h00;
		ram[15'h663] =  8'h00;
		ram[15'h664] =  8'h00;
		ram[15'h665] =  8'h00;
		ram[15'h666] =  8'h00;
		ram[15'h667] =  8'h00;
		ram[15'h668] =  8'h00;
		ram[15'h669] =  8'h00;
		ram[15'h66A] =  8'h00;
		ram[15'h66B] =  8'h00;
		ram[15'h66C] =  8'h00;
		ram[15'h66D] =  8'h00;
		ram[15'h66E] =  8'h00;
		ram[15'h66F] =  8'h00;
		ram[15'h670] =  8'h00;
		ram[15'h671] =  8'h00;
		ram[15'h672] =  8'h00;
		ram[15'h673] =  8'hD7;
		ram[15'h674] =  8'h00;
		ram[15'h675] =  8'h00;
		ram[15'h676] =  8'h00;
		ram[15'h677] =  8'h5F;
		ram[15'h678] =  8'h68;
		ram[15'h679] =  8'h22;
		ram[15'h67A] =  8'h64;
		ram[15'h67B] =  8'h3C;
		ram[15'h67C] =  8'h69;
		ram[15'h67D] =  8'h6E;
		ram[15'h67E] =  8'h63;
		ram[15'h67F] =  8'h2C;
		ram[15'h680] =  8'h64;
		ram[15'h681] =  8'h65;
		ram[15'h682] =  8'h63;
		ram[15'h683] =  8'h3E;
		ram[15'h684] =  8'h20;
		ram[15'h685] =  8'h62;
		ram[15'h686] =  8'h2E;
		ram[15'h687] =  8'h2E;
		ram[15'h688] =  8'h2E;
		ram[15'h689] =  8'h2E;
		ram[15'h68A] =  8'h2E;
		ram[15'h68B] =  8'h2E;
		ram[15'h68C] =  8'h2E;
		ram[15'h68D] =  8'h2E;
		ram[15'h68E] =  8'h2E;
		ram[15'h68F] =  8'h2E;
		ram[15'h690] =  8'h2E;
		ram[15'h691] =  8'h2E;
		ram[15'h692] =  8'h2E;
		ram[15'h693] =  8'h2E;
		ram[15'h694] =  8'h2E;
		ram[15'h695] =  8'h2E;
		ram[15'h696] =  8'h2E;
		ram[15'h697] =  8'h2E;
		ram[15'h698] =  8'h2E;
		ram[15'h699] =  8'h24;
		ram[15'h69A] =  8'hD7;
		ram[15'h69B] =  8'h03;
		ram[15'h69C] =  8'h00;
		ram[15'h69D] =  8'h00;
		ram[15'h69E] =  8'h00;
		ram[15'h69F] =  8'h97;
		ram[15'h6A0] =  8'hCD;
		ram[15'h6A1] =  8'hAB;
		ram[15'h6A2] =  8'h44;
		ram[15'h6A3] =  8'hC9;
		ram[15'h6A4] =  8'h8D;
		ram[15'h6A5] =  8'hE3;
		ram[15'h6A6] =  8'hE3;
		ram[15'h6A7] =  8'hCC;
		ram[15'h6A8] =  8'h11;
		ram[15'h6A9] =  8'hA4;
		ram[15'h6AA] =  8'hE8;
		ram[15'h6AB] =  8'h02;
		ram[15'h6AC] =  8'h49;
		ram[15'h6AD] =  8'h4D;
		ram[15'h6AE] =  8'h2A;
		ram[15'h6AF] =  8'h08;
		ram[15'h6B0] =  8'h00;
		ram[15'h6B1] =  8'h00;
		ram[15'h6B2] =  8'h00;
		ram[15'h6B3] =  8'h00;
		ram[15'h6B4] =  8'h00;
		ram[15'h6B5] =  8'h00;
		ram[15'h6B6] =  8'h00;
		ram[15'h6B7] =  8'h00;
		ram[15'h6B8] =  8'h00;
		ram[15'h6B9] =  8'h00;
		ram[15'h6BA] =  8'h00;
		ram[15'h6BB] =  8'h00;
		ram[15'h6BC] =  8'h00;
		ram[15'h6BD] =  8'h21;
		ram[15'h6BE] =  8'hF8;
		ram[15'h6BF] =  8'h00;
		ram[15'h6C0] =  8'h00;
		ram[15'h6C1] =  8'h00;
		ram[15'h6C2] =  8'h00;
		ram[15'h6C3] =  8'h00;
		ram[15'h6C4] =  8'h00;
		ram[15'h6C5] =  8'h00;
		ram[15'h6C6] =  8'h00;
		ram[15'h6C7] =  8'h00;
		ram[15'h6C8] =  8'h00;
		ram[15'h6C9] =  8'h00;
		ram[15'h6CA] =  8'h00;
		ram[15'h6CB] =  8'h00;
		ram[15'h6CC] =  8'h00;
		ram[15'h6CD] =  8'h00;
		ram[15'h6CE] =  8'h00;
		ram[15'h6CF] =  8'h00;
		ram[15'h6D0] =  8'h00;
		ram[15'h6D1] =  8'h00;
		ram[15'h6D2] =  8'h00;
		ram[15'h6D3] =  8'hD7;
		ram[15'h6D4] =  8'h00;
		ram[15'h6D5] =  8'h00;
		ram[15'h6D6] =  8'h00;
		ram[15'h6D7] =  8'hD2;
		ram[15'h6D8] =  8'hAE;
		ram[15'h6D9] =  8'h3B;
		ram[15'h6DA] =  8'hEC;
		ram[15'h6DB] =  8'h3C;
		ram[15'h6DC] =  8'h69;
		ram[15'h6DD] =  8'h6E;
		ram[15'h6DE] =  8'h63;
		ram[15'h6DF] =  8'h2C;
		ram[15'h6E0] =  8'h64;
		ram[15'h6E1] =  8'h65;
		ram[15'h6E2] =  8'h63;
		ram[15'h6E3] =  8'h3E;
		ram[15'h6E4] =  8'h20;
		ram[15'h6E5] =  8'h62;
		ram[15'h6E6] =  8'h63;
		ram[15'h6E7] =  8'h2E;
		ram[15'h6E8] =  8'h2E;
		ram[15'h6E9] =  8'h2E;
		ram[15'h6EA] =  8'h2E;
		ram[15'h6EB] =  8'h2E;
		ram[15'h6EC] =  8'h2E;
		ram[15'h6ED] =  8'h2E;
		ram[15'h6EE] =  8'h2E;
		ram[15'h6EF] =  8'h2E;
		ram[15'h6F0] =  8'h2E;
		ram[15'h6F1] =  8'h2E;
		ram[15'h6F2] =  8'h2E;
		ram[15'h6F3] =  8'h2E;
		ram[15'h6F4] =  8'h2E;
		ram[15'h6F5] =  8'h2E;
		ram[15'h6F6] =  8'h2E;
		ram[15'h6F7] =  8'h2E;
		ram[15'h6F8] =  8'h2E;
		ram[15'h6F9] =  8'h24;
		ram[15'h6FA] =  8'hD7;
		ram[15'h6FB] =  8'h0C;
		ram[15'h6FC] =  8'h00;
		ram[15'h6FD] =  8'h00;
		ram[15'h6FE] =  8'h00;
		ram[15'h6FF] =  8'h89;
		ram[15'h700] =  8'hD7;
		ram[15'h701] =  8'h35;
		ram[15'h702] =  8'h09;
		ram[15'h703] =  8'h5B;
		ram[15'h704] =  8'h05;
		ram[15'h705] =  8'h85;
		ram[15'h706] =  8'h9F;
		ram[15'h707] =  8'h27;
		ram[15'h708] =  8'h8B;
		ram[15'h709] =  8'h08;
		ram[15'h70A] =  8'hD2;
		ram[15'h70B] =  8'h95;
		ram[15'h70C] =  8'h05;
		ram[15'h70D] =  8'h60;
		ram[15'h70E] =  8'h06;
		ram[15'h70F] =  8'h01;
		ram[15'h710] =  8'h00;
		ram[15'h711] =  8'h00;
		ram[15'h712] =  8'h00;
		ram[15'h713] =  8'h00;
		ram[15'h714] =  8'h00;
		ram[15'h715] =  8'h00;
		ram[15'h716] =  8'h00;
		ram[15'h717] =  8'h00;
		ram[15'h718] =  8'h00;
		ram[15'h719] =  8'h00;
		ram[15'h71A] =  8'h00;
		ram[15'h71B] =  8'h00;
		ram[15'h71C] =  8'h00;
		ram[15'h71D] =  8'hFF;
		ram[15'h71E] =  8'h00;
		ram[15'h71F] =  8'h00;
		ram[15'h720] =  8'h00;
		ram[15'h721] =  8'h00;
		ram[15'h722] =  8'h00;
		ram[15'h723] =  8'h00;
		ram[15'h724] =  8'h00;
		ram[15'h725] =  8'h00;
		ram[15'h726] =  8'h00;
		ram[15'h727] =  8'h00;
		ram[15'h728] =  8'h00;
		ram[15'h729] =  8'h00;
		ram[15'h72A] =  8'h00;
		ram[15'h72B] =  8'h00;
		ram[15'h72C] =  8'h00;
		ram[15'h72D] =  8'h00;
		ram[15'h72E] =  8'h00;
		ram[15'h72F] =  8'h00;
		ram[15'h730] =  8'h00;
		ram[15'h731] =  8'h00;
		ram[15'h732] =  8'h00;
		ram[15'h733] =  8'hD7;
		ram[15'h734] =  8'h00;
		ram[15'h735] =  8'h00;
		ram[15'h736] =  8'h00;
		ram[15'h737] =  8'hC2;
		ram[15'h738] =  8'h84;
		ram[15'h739] =  8'h55;
		ram[15'h73A] =  8'h4C;
		ram[15'h73B] =  8'h3C;
		ram[15'h73C] =  8'h69;
		ram[15'h73D] =  8'h6E;
		ram[15'h73E] =  8'h63;
		ram[15'h73F] =  8'h2C;
		ram[15'h740] =  8'h64;
		ram[15'h741] =  8'h65;
		ram[15'h742] =  8'h63;
		ram[15'h743] =  8'h3E;
		ram[15'h744] =  8'h20;
		ram[15'h745] =  8'h63;
		ram[15'h746] =  8'h2E;
		ram[15'h747] =  8'h2E;
		ram[15'h748] =  8'h2E;
		ram[15'h749] =  8'h2E;
		ram[15'h74A] =  8'h2E;
		ram[15'h74B] =  8'h2E;
		ram[15'h74C] =  8'h2E;
		ram[15'h74D] =  8'h2E;
		ram[15'h74E] =  8'h2E;
		ram[15'h74F] =  8'h2E;
		ram[15'h750] =  8'h2E;
		ram[15'h751] =  8'h2E;
		ram[15'h752] =  8'h2E;
		ram[15'h753] =  8'h2E;
		ram[15'h754] =  8'h2E;
		ram[15'h755] =  8'h2E;
		ram[15'h756] =  8'h2E;
		ram[15'h757] =  8'h2E;
		ram[15'h758] =  8'h2E;
		ram[15'h759] =  8'h24;
		ram[15'h75A] =  8'hD7;
		ram[15'h75B] =  8'h14;
		ram[15'h75C] =  8'h00;
		ram[15'h75D] =  8'h00;
		ram[15'h75E] =  8'h00;
		ram[15'h75F] =  8'hEA;
		ram[15'h760] =  8'hA0;
		ram[15'h761] =  8'hBA;
		ram[15'h762] =  8'h5F;
		ram[15'h763] =  8'hFB;
		ram[15'h764] =  8'h65;
		ram[15'h765] =  8'h1C;
		ram[15'h766] =  8'h98;
		ram[15'h767] =  8'hCC;
		ram[15'h768] =  8'h38;
		ram[15'h769] =  8'hBC;
		ram[15'h76A] =  8'hDE;
		ram[15'h76B] =  8'h43;
		ram[15'h76C] =  8'h5C;
		ram[15'h76D] =  8'hBD;
		ram[15'h76E] =  8'h03;
		ram[15'h76F] =  8'h01;
		ram[15'h770] =  8'h00;
		ram[15'h771] =  8'h00;
		ram[15'h772] =  8'h00;
		ram[15'h773] =  8'h00;
		ram[15'h774] =  8'h00;
		ram[15'h775] =  8'h00;
		ram[15'h776] =  8'h00;
		ram[15'h777] =  8'h00;
		ram[15'h778] =  8'h00;
		ram[15'h779] =  8'h00;
		ram[15'h77A] =  8'h00;
		ram[15'h77B] =  8'h00;
		ram[15'h77C] =  8'hFF;
		ram[15'h77D] =  8'h00;
		ram[15'h77E] =  8'h00;
		ram[15'h77F] =  8'h00;
		ram[15'h780] =  8'h00;
		ram[15'h781] =  8'h00;
		ram[15'h782] =  8'h00;
		ram[15'h783] =  8'h00;
		ram[15'h784] =  8'h00;
		ram[15'h785] =  8'h00;
		ram[15'h786] =  8'h00;
		ram[15'h787] =  8'h00;
		ram[15'h788] =  8'h00;
		ram[15'h789] =  8'h00;
		ram[15'h78A] =  8'h00;
		ram[15'h78B] =  8'h00;
		ram[15'h78C] =  8'h00;
		ram[15'h78D] =  8'h00;
		ram[15'h78E] =  8'h00;
		ram[15'h78F] =  8'h00;
		ram[15'h790] =  8'h00;
		ram[15'h791] =  8'h00;
		ram[15'h792] =  8'h00;
		ram[15'h793] =  8'hD7;
		ram[15'h794] =  8'h00;
		ram[15'h795] =  8'h00;
		ram[15'h796] =  8'h00;
		ram[15'h797] =  8'h45;
		ram[15'h798] =  8'h23;
		ram[15'h799] =  8'hDE;
		ram[15'h79A] =  8'h10;
		ram[15'h79B] =  8'h3C;
		ram[15'h79C] =  8'h69;
		ram[15'h79D] =  8'h6E;
		ram[15'h79E] =  8'h63;
		ram[15'h79F] =  8'h2C;
		ram[15'h7A0] =  8'h64;
		ram[15'h7A1] =  8'h65;
		ram[15'h7A2] =  8'h63;
		ram[15'h7A3] =  8'h3E;
		ram[15'h7A4] =  8'h20;
		ram[15'h7A5] =  8'h64;
		ram[15'h7A6] =  8'h2E;
		ram[15'h7A7] =  8'h2E;
		ram[15'h7A8] =  8'h2E;
		ram[15'h7A9] =  8'h2E;
		ram[15'h7AA] =  8'h2E;
		ram[15'h7AB] =  8'h2E;
		ram[15'h7AC] =  8'h2E;
		ram[15'h7AD] =  8'h2E;
		ram[15'h7AE] =  8'h2E;
		ram[15'h7AF] =  8'h2E;
		ram[15'h7B0] =  8'h2E;
		ram[15'h7B1] =  8'h2E;
		ram[15'h7B2] =  8'h2E;
		ram[15'h7B3] =  8'h2E;
		ram[15'h7B4] =  8'h2E;
		ram[15'h7B5] =  8'h2E;
		ram[15'h7B6] =  8'h2E;
		ram[15'h7B7] =  8'h2E;
		ram[15'h7B8] =  8'h2E;
		ram[15'h7B9] =  8'h24;
		ram[15'h7BA] =  8'hD7;
		ram[15'h7BB] =  8'h13;
		ram[15'h7BC] =  8'h00;
		ram[15'h7BD] =  8'h00;
		ram[15'h7BE] =  8'h00;
		ram[15'h7BF] =  8'h2E;
		ram[15'h7C0] =  8'h34;
		ram[15'h7C1] =  8'h1D;
		ram[15'h7C2] =  8'h13;
		ram[15'h7C3] =  8'hC9;
		ram[15'h7C4] =  8'h28;
		ram[15'h7C5] =  8'hCA;
		ram[15'h7C6] =  8'h0A;
		ram[15'h7C7] =  8'h67;
		ram[15'h7C8] =  8'h99;
		ram[15'h7C9] =  8'h2E;
		ram[15'h7CA] =  8'h3A;
		ram[15'h7CB] =  8'h92;
		ram[15'h7CC] =  8'hF6;
		ram[15'h7CD] =  8'h54;
		ram[15'h7CE] =  8'h9D;
		ram[15'h7CF] =  8'h08;
		ram[15'h7D0] =  8'h00;
		ram[15'h7D1] =  8'h00;
		ram[15'h7D2] =  8'h00;
		ram[15'h7D3] =  8'h00;
		ram[15'h7D4] =  8'h00;
		ram[15'h7D5] =  8'h00;
		ram[15'h7D6] =  8'h00;
		ram[15'h7D7] =  8'h00;
		ram[15'h7D8] =  8'h00;
		ram[15'h7D9] =  8'h00;
		ram[15'h7DA] =  8'h00;
		ram[15'h7DB] =  8'h21;
		ram[15'h7DC] =  8'hF8;
		ram[15'h7DD] =  8'h00;
		ram[15'h7DE] =  8'h00;
		ram[15'h7DF] =  8'h00;
		ram[15'h7E0] =  8'h00;
		ram[15'h7E1] =  8'h00;
		ram[15'h7E2] =  8'h00;
		ram[15'h7E3] =  8'h00;
		ram[15'h7E4] =  8'h00;
		ram[15'h7E5] =  8'h00;
		ram[15'h7E6] =  8'h00;
		ram[15'h7E7] =  8'h00;
		ram[15'h7E8] =  8'h00;
		ram[15'h7E9] =  8'h00;
		ram[15'h7EA] =  8'h00;
		ram[15'h7EB] =  8'h00;
		ram[15'h7EC] =  8'h00;
		ram[15'h7ED] =  8'h00;
		ram[15'h7EE] =  8'h00;
		ram[15'h7EF] =  8'h00;
		ram[15'h7F0] =  8'h00;
		ram[15'h7F1] =  8'h00;
		ram[15'h7F2] =  8'h00;
		ram[15'h7F3] =  8'hD7;
		ram[15'h7F4] =  8'h00;
		ram[15'h7F5] =  8'h00;
		ram[15'h7F6] =  8'h00;
		ram[15'h7F7] =  8'hAE;
		ram[15'h7F8] =  8'hC6;
		ram[15'h7F9] =  8'hD4;
		ram[15'h7FA] =  8'h2C;
		ram[15'h7FB] =  8'h3C;
		ram[15'h7FC] =  8'h69;
		ram[15'h7FD] =  8'h6E;
		ram[15'h7FE] =  8'h63;
		ram[15'h7FF] =  8'h2C;
		ram[15'h800] =  8'h64;
		ram[15'h801] =  8'h65;
		ram[15'h802] =  8'h63;
		ram[15'h803] =  8'h3E;
		ram[15'h804] =  8'h20;
		ram[15'h805] =  8'h64;
		ram[15'h806] =  8'h65;
		ram[15'h807] =  8'h2E;
		ram[15'h808] =  8'h2E;
		ram[15'h809] =  8'h2E;
		ram[15'h80A] =  8'h2E;
		ram[15'h80B] =  8'h2E;
		ram[15'h80C] =  8'h2E;
		ram[15'h80D] =  8'h2E;
		ram[15'h80E] =  8'h2E;
		ram[15'h80F] =  8'h2E;
		ram[15'h810] =  8'h2E;
		ram[15'h811] =  8'h2E;
		ram[15'h812] =  8'h2E;
		ram[15'h813] =  8'h2E;
		ram[15'h814] =  8'h2E;
		ram[15'h815] =  8'h2E;
		ram[15'h816] =  8'h2E;
		ram[15'h817] =  8'h2E;
		ram[15'h818] =  8'h2E;
		ram[15'h819] =  8'h24;
		ram[15'h81A] =  8'hD7;
		ram[15'h81B] =  8'h1C;
		ram[15'h81C] =  8'h00;
		ram[15'h81D] =  8'h00;
		ram[15'h81E] =  8'h00;
		ram[15'h81F] =  8'h2F;
		ram[15'h820] =  8'h60;
		ram[15'h821] =  8'h0D;
		ram[15'h822] =  8'h4C;
		ram[15'h823] =  8'h02;
		ram[15'h824] =  8'h24;
		ram[15'h825] =  8'hF5;
		ram[15'h826] =  8'hE2;
		ram[15'h827] =  8'hF4;
		ram[15'h828] =  8'hA0;
		ram[15'h829] =  8'h0A;
		ram[15'h82A] =  8'hA1;
		ram[15'h82B] =  8'h13;
		ram[15'h82C] =  8'h32;
		ram[15'h82D] =  8'h25;
		ram[15'h82E] =  8'h59;
		ram[15'h82F] =  8'h01;
		ram[15'h830] =  8'h00;
		ram[15'h831] =  8'h00;
		ram[15'h832] =  8'h00;
		ram[15'h833] =  8'h00;
		ram[15'h834] =  8'h00;
		ram[15'h835] =  8'h00;
		ram[15'h836] =  8'h00;
		ram[15'h837] =  8'h00;
		ram[15'h838] =  8'h00;
		ram[15'h839] =  8'h00;
		ram[15'h83A] =  8'h00;
		ram[15'h83B] =  8'hFF;
		ram[15'h83C] =  8'h00;
		ram[15'h83D] =  8'h00;
		ram[15'h83E] =  8'h00;
		ram[15'h83F] =  8'h00;
		ram[15'h840] =  8'h00;
		ram[15'h841] =  8'h00;
		ram[15'h842] =  8'h00;
		ram[15'h843] =  8'h00;
		ram[15'h844] =  8'h00;
		ram[15'h845] =  8'h00;
		ram[15'h846] =  8'h00;
		ram[15'h847] =  8'h00;
		ram[15'h848] =  8'h00;
		ram[15'h849] =  8'h00;
		ram[15'h84A] =  8'h00;
		ram[15'h84B] =  8'h00;
		ram[15'h84C] =  8'h00;
		ram[15'h84D] =  8'h00;
		ram[15'h84E] =  8'h00;
		ram[15'h84F] =  8'h00;
		ram[15'h850] =  8'h00;
		ram[15'h851] =  8'h00;
		ram[15'h852] =  8'h00;
		ram[15'h853] =  8'hD7;
		ram[15'h854] =  8'h00;
		ram[15'h855] =  8'h00;
		ram[15'h856] =  8'h00;
		ram[15'h857] =  8'hE1;
		ram[15'h858] =  8'h75;
		ram[15'h859] =  8'hAF;
		ram[15'h85A] =  8'hCC;
		ram[15'h85B] =  8'h3C;
		ram[15'h85C] =  8'h69;
		ram[15'h85D] =  8'h6E;
		ram[15'h85E] =  8'h63;
		ram[15'h85F] =  8'h2C;
		ram[15'h860] =  8'h64;
		ram[15'h861] =  8'h65;
		ram[15'h862] =  8'h63;
		ram[15'h863] =  8'h3E;
		ram[15'h864] =  8'h20;
		ram[15'h865] =  8'h65;
		ram[15'h866] =  8'h2E;
		ram[15'h867] =  8'h2E;
		ram[15'h868] =  8'h2E;
		ram[15'h869] =  8'h2E;
		ram[15'h86A] =  8'h2E;
		ram[15'h86B] =  8'h2E;
		ram[15'h86C] =  8'h2E;
		ram[15'h86D] =  8'h2E;
		ram[15'h86E] =  8'h2E;
		ram[15'h86F] =  8'h2E;
		ram[15'h870] =  8'h2E;
		ram[15'h871] =  8'h2E;
		ram[15'h872] =  8'h2E;
		ram[15'h873] =  8'h2E;
		ram[15'h874] =  8'h2E;
		ram[15'h875] =  8'h2E;
		ram[15'h876] =  8'h2E;
		ram[15'h877] =  8'h2E;
		ram[15'h878] =  8'h2E;
		ram[15'h879] =  8'h24;
		ram[15'h87A] =  8'hD7;
		ram[15'h87B] =  8'h24;
		ram[15'h87C] =  8'h00;
		ram[15'h87D] =  8'h00;
		ram[15'h87E] =  8'h00;
		ram[15'h87F] =  8'h06;
		ram[15'h880] =  8'h15;
		ram[15'h881] =  8'hEB;
		ram[15'h882] =  8'hF2;
		ram[15'h883] =  8'hDD;
		ram[15'h884] =  8'hE8;
		ram[15'h885] =  8'h2B;
		ram[15'h886] =  8'h26;
		ram[15'h887] =  8'hA6;
		ram[15'h888] =  8'h11;
		ram[15'h889] =  8'h1A;
		ram[15'h88A] =  8'hBC;
		ram[15'h88B] =  8'h17;
		ram[15'h88C] =  8'h06;
		ram[15'h88D] =  8'h18;
		ram[15'h88E] =  8'h28;
		ram[15'h88F] =  8'h01;
		ram[15'h890] =  8'h00;
		ram[15'h891] =  8'h00;
		ram[15'h892] =  8'h00;
		ram[15'h893] =  8'h00;
		ram[15'h894] =  8'h00;
		ram[15'h895] =  8'h00;
		ram[15'h896] =  8'h00;
		ram[15'h897] =  8'h00;
		ram[15'h898] =  8'h00;
		ram[15'h899] =  8'h00;
		ram[15'h89A] =  8'hFF;
		ram[15'h89B] =  8'h00;
		ram[15'h89C] =  8'h00;
		ram[15'h89D] =  8'h00;
		ram[15'h89E] =  8'h00;
		ram[15'h89F] =  8'h00;
		ram[15'h8A0] =  8'h00;
		ram[15'h8A1] =  8'h00;
		ram[15'h8A2] =  8'h00;
		ram[15'h8A3] =  8'h00;
		ram[15'h8A4] =  8'h00;
		ram[15'h8A5] =  8'h00;
		ram[15'h8A6] =  8'h00;
		ram[15'h8A7] =  8'h00;
		ram[15'h8A8] =  8'h00;
		ram[15'h8A9] =  8'h00;
		ram[15'h8AA] =  8'h00;
		ram[15'h8AB] =  8'h00;
		ram[15'h8AC] =  8'h00;
		ram[15'h8AD] =  8'h00;
		ram[15'h8AE] =  8'h00;
		ram[15'h8AF] =  8'h00;
		ram[15'h8B0] =  8'h00;
		ram[15'h8B1] =  8'h00;
		ram[15'h8B2] =  8'h00;
		ram[15'h8B3] =  8'hD7;
		ram[15'h8B4] =  8'h00;
		ram[15'h8B5] =  8'h00;
		ram[15'h8B6] =  8'h00;
		ram[15'h8B7] =  8'h1C;
		ram[15'h8B8] =  8'hED;
		ram[15'h8B9] =  8'h84;
		ram[15'h8BA] =  8'h7D;
		ram[15'h8BB] =  8'h3C;
		ram[15'h8BC] =  8'h69;
		ram[15'h8BD] =  8'h6E;
		ram[15'h8BE] =  8'h63;
		ram[15'h8BF] =  8'h2C;
		ram[15'h8C0] =  8'h64;
		ram[15'h8C1] =  8'h65;
		ram[15'h8C2] =  8'h63;
		ram[15'h8C3] =  8'h3E;
		ram[15'h8C4] =  8'h20;
		ram[15'h8C5] =  8'h68;
		ram[15'h8C6] =  8'h2E;
		ram[15'h8C7] =  8'h2E;
		ram[15'h8C8] =  8'h2E;
		ram[15'h8C9] =  8'h2E;
		ram[15'h8CA] =  8'h2E;
		ram[15'h8CB] =  8'h2E;
		ram[15'h8CC] =  8'h2E;
		ram[15'h8CD] =  8'h2E;
		ram[15'h8CE] =  8'h2E;
		ram[15'h8CF] =  8'h2E;
		ram[15'h8D0] =  8'h2E;
		ram[15'h8D1] =  8'h2E;
		ram[15'h8D2] =  8'h2E;
		ram[15'h8D3] =  8'h2E;
		ram[15'h8D4] =  8'h2E;
		ram[15'h8D5] =  8'h2E;
		ram[15'h8D6] =  8'h2E;
		ram[15'h8D7] =  8'h2E;
		ram[15'h8D8] =  8'h2E;
		ram[15'h8D9] =  8'h24;
		ram[15'h8DA] =  8'hD7;
		ram[15'h8DB] =  8'h23;
		ram[15'h8DC] =  8'h00;
		ram[15'h8DD] =  8'h00;
		ram[15'h8DE] =  8'h00;
		ram[15'h8DF] =  8'hF4;
		ram[15'h8E0] =  8'hC3;
		ram[15'h8E1] =  8'hA5;
		ram[15'h8E2] =  8'h07;
		ram[15'h8E3] =  8'h6D;
		ram[15'h8E4] =  8'h1B;
		ram[15'h8E5] =  8'h04;
		ram[15'h8E6] =  8'h4F;
		ram[15'h8E7] =  8'hC2;
		ram[15'h8E8] =  8'hE2;
		ram[15'h8E9] =  8'h2A;
		ram[15'h8EA] =  8'h82;
		ram[15'h8EB] =  8'h57;
		ram[15'h8EC] =  8'hE0;
		ram[15'h8ED] =  8'hE1;
		ram[15'h8EE] =  8'hC3;
		ram[15'h8EF] =  8'h08;
		ram[15'h8F0] =  8'h00;
		ram[15'h8F1] =  8'h00;
		ram[15'h8F2] =  8'h00;
		ram[15'h8F3] =  8'h00;
		ram[15'h8F4] =  8'h00;
		ram[15'h8F5] =  8'h00;
		ram[15'h8F6] =  8'h00;
		ram[15'h8F7] =  8'h00;
		ram[15'h8F8] =  8'h00;
		ram[15'h8F9] =  8'h21;
		ram[15'h8FA] =  8'hF8;
		ram[15'h8FB] =  8'h00;
		ram[15'h8FC] =  8'h00;
		ram[15'h8FD] =  8'h00;
		ram[15'h8FE] =  8'h00;
		ram[15'h8FF] =  8'h00;
		ram[15'h900] =  8'h00;
		ram[15'h901] =  8'h00;
		ram[15'h902] =  8'h00;
		ram[15'h903] =  8'h00;
		ram[15'h904] =  8'h00;
		ram[15'h905] =  8'h00;
		ram[15'h906] =  8'h00;
		ram[15'h907] =  8'h00;
		ram[15'h908] =  8'h00;
		ram[15'h909] =  8'h00;
		ram[15'h90A] =  8'h00;
		ram[15'h90B] =  8'h00;
		ram[15'h90C] =  8'h00;
		ram[15'h90D] =  8'h00;
		ram[15'h90E] =  8'h00;
		ram[15'h90F] =  8'h00;
		ram[15'h910] =  8'h00;
		ram[15'h911] =  8'h00;
		ram[15'h912] =  8'h00;
		ram[15'h913] =  8'hD7;
		ram[15'h914] =  8'h00;
		ram[15'h915] =  8'h00;
		ram[15'h916] =  8'h00;
		ram[15'h917] =  8'hFC;
		ram[15'h918] =  8'h0D;
		ram[15'h919] =  8'h6D;
		ram[15'h91A] =  8'h4A;
		ram[15'h91B] =  8'h3C;
		ram[15'h91C] =  8'h69;
		ram[15'h91D] =  8'h6E;
		ram[15'h91E] =  8'h63;
		ram[15'h91F] =  8'h2C;
		ram[15'h920] =  8'h64;
		ram[15'h921] =  8'h65;
		ram[15'h922] =  8'h63;
		ram[15'h923] =  8'h3E;
		ram[15'h924] =  8'h20;
		ram[15'h925] =  8'h68;
		ram[15'h926] =  8'h6C;
		ram[15'h927] =  8'h2E;
		ram[15'h928] =  8'h2E;
		ram[15'h929] =  8'h2E;
		ram[15'h92A] =  8'h2E;
		ram[15'h92B] =  8'h2E;
		ram[15'h92C] =  8'h2E;
		ram[15'h92D] =  8'h2E;
		ram[15'h92E] =  8'h2E;
		ram[15'h92F] =  8'h2E;
		ram[15'h930] =  8'h2E;
		ram[15'h931] =  8'h2E;
		ram[15'h932] =  8'h2E;
		ram[15'h933] =  8'h2E;
		ram[15'h934] =  8'h2E;
		ram[15'h935] =  8'h2E;
		ram[15'h936] =  8'h2E;
		ram[15'h937] =  8'h2E;
		ram[15'h938] =  8'h2E;
		ram[15'h939] =  8'h24;
		ram[15'h93A] =  8'hD7;
		ram[15'h93B] =  8'hDD;
		ram[15'h93C] =  8'h23;
		ram[15'h93D] =  8'h00;
		ram[15'h93E] =  8'h00;
		ram[15'h93F] =  8'h3C;
		ram[15'h940] =  8'hBC;
		ram[15'h941] =  8'h9B;
		ram[15'h942] =  8'h0D;
		ram[15'h943] =  8'h81;
		ram[15'h944] =  8'hE0;
		ram[15'h945] =  8'hFD;
		ram[15'h946] =  8'hAD;
		ram[15'h947] =  8'h7F;
		ram[15'h948] =  8'h9A;
		ram[15'h949] =  8'hE5;
		ram[15'h94A] =  8'h96;
		ram[15'h94B] =  8'h13;
		ram[15'h94C] =  8'h85;
		ram[15'h94D] =  8'hE2;
		ram[15'h94E] =  8'h0B;
		ram[15'h94F] =  8'h00;
		ram[15'h950] =  8'h08;
		ram[15'h951] =  8'h00;
		ram[15'h952] =  8'h00;
		ram[15'h953] =  8'h00;
		ram[15'h954] =  8'h00;
		ram[15'h955] =  8'h00;
		ram[15'h956] =  8'h00;
		ram[15'h957] =  8'h21;
		ram[15'h958] =  8'hF8;
		ram[15'h959] =  8'h00;
		ram[15'h95A] =  8'h00;
		ram[15'h95B] =  8'h00;
		ram[15'h95C] =  8'h00;
		ram[15'h95D] =  8'h00;
		ram[15'h95E] =  8'h00;
		ram[15'h95F] =  8'h00;
		ram[15'h960] =  8'h00;
		ram[15'h961] =  8'h00;
		ram[15'h962] =  8'h00;
		ram[15'h963] =  8'h00;
		ram[15'h964] =  8'h00;
		ram[15'h965] =  8'h00;
		ram[15'h966] =  8'h00;
		ram[15'h967] =  8'h00;
		ram[15'h968] =  8'h00;
		ram[15'h969] =  8'h00;
		ram[15'h96A] =  8'h00;
		ram[15'h96B] =  8'h00;
		ram[15'h96C] =  8'h00;
		ram[15'h96D] =  8'h00;
		ram[15'h96E] =  8'h00;
		ram[15'h96F] =  8'h00;
		ram[15'h970] =  8'h00;
		ram[15'h971] =  8'h00;
		ram[15'h972] =  8'h00;
		ram[15'h973] =  8'hD7;
		ram[15'h974] =  8'h00;
		ram[15'h975] =  8'h00;
		ram[15'h976] =  8'h00;
		ram[15'h977] =  8'hA5;
		ram[15'h978] =  8'h4D;
		ram[15'h979] =  8'hBE;
		ram[15'h97A] =  8'h31;
		ram[15'h97B] =  8'h3C;
		ram[15'h97C] =  8'h69;
		ram[15'h97D] =  8'h6E;
		ram[15'h97E] =  8'h63;
		ram[15'h97F] =  8'h2C;
		ram[15'h980] =  8'h64;
		ram[15'h981] =  8'h65;
		ram[15'h982] =  8'h63;
		ram[15'h983] =  8'h3E;
		ram[15'h984] =  8'h20;
		ram[15'h985] =  8'h69;
		ram[15'h986] =  8'h78;
		ram[15'h987] =  8'h2E;
		ram[15'h988] =  8'h2E;
		ram[15'h989] =  8'h2E;
		ram[15'h98A] =  8'h2E;
		ram[15'h98B] =  8'h2E;
		ram[15'h98C] =  8'h2E;
		ram[15'h98D] =  8'h2E;
		ram[15'h98E] =  8'h2E;
		ram[15'h98F] =  8'h2E;
		ram[15'h990] =  8'h2E;
		ram[15'h991] =  8'h2E;
		ram[15'h992] =  8'h2E;
		ram[15'h993] =  8'h2E;
		ram[15'h994] =  8'h2E;
		ram[15'h995] =  8'h2E;
		ram[15'h996] =  8'h2E;
		ram[15'h997] =  8'h2E;
		ram[15'h998] =  8'h2E;
		ram[15'h999] =  8'h24;
		ram[15'h99A] =  8'hD7;
		ram[15'h99B] =  8'hFD;
		ram[15'h99C] =  8'h23;
		ram[15'h99D] =  8'h00;
		ram[15'h99E] =  8'h00;
		ram[15'h99F] =  8'h02;
		ram[15'h9A0] =  8'h94;
		ram[15'h9A1] =  8'h7A;
		ram[15'h9A2] =  8'h63;
		ram[15'h9A3] =  8'h82;
		ram[15'h9A4] =  8'h31;
		ram[15'h9A5] =  8'h5A;
		ram[15'h9A6] =  8'hC6;
		ram[15'h9A7] =  8'hE9;
		ram[15'h9A8] =  8'hB2;
		ram[15'h9A9] =  8'hB4;
		ram[15'h9AA] =  8'hAB;
		ram[15'h9AB] =  8'h16;
		ram[15'h9AC] =  8'hF2;
		ram[15'h9AD] =  8'h05;
		ram[15'h9AE] =  8'h6D;
		ram[15'h9AF] =  8'h00;
		ram[15'h9B0] =  8'h08;
		ram[15'h9B1] =  8'h00;
		ram[15'h9B2] =  8'h00;
		ram[15'h9B3] =  8'h00;
		ram[15'h9B4] =  8'h00;
		ram[15'h9B5] =  8'h21;
		ram[15'h9B6] =  8'hF8;
		ram[15'h9B7] =  8'h00;
		ram[15'h9B8] =  8'h00;
		ram[15'h9B9] =  8'h00;
		ram[15'h9BA] =  8'h00;
		ram[15'h9BB] =  8'h00;
		ram[15'h9BC] =  8'h00;
		ram[15'h9BD] =  8'h00;
		ram[15'h9BE] =  8'h00;
		ram[15'h9BF] =  8'h00;
		ram[15'h9C0] =  8'h00;
		ram[15'h9C1] =  8'h00;
		ram[15'h9C2] =  8'h00;
		ram[15'h9C3] =  8'h00;
		ram[15'h9C4] =  8'h00;
		ram[15'h9C5] =  8'h00;
		ram[15'h9C6] =  8'h00;
		ram[15'h9C7] =  8'h00;
		ram[15'h9C8] =  8'h00;
		ram[15'h9C9] =  8'h00;
		ram[15'h9CA] =  8'h00;
		ram[15'h9CB] =  8'h00;
		ram[15'h9CC] =  8'h00;
		ram[15'h9CD] =  8'h00;
		ram[15'h9CE] =  8'h00;
		ram[15'h9CF] =  8'h00;
		ram[15'h9D0] =  8'h00;
		ram[15'h9D1] =  8'h00;
		ram[15'h9D2] =  8'h00;
		ram[15'h9D3] =  8'hD7;
		ram[15'h9D4] =  8'h00;
		ram[15'h9D5] =  8'h00;
		ram[15'h9D6] =  8'h00;
		ram[15'h9D7] =  8'h50;
		ram[15'h9D8] =  8'h5D;
		ram[15'h9D9] =  8'h51;
		ram[15'h9DA] =  8'hA3;
		ram[15'h9DB] =  8'h3C;
		ram[15'h9DC] =  8'h69;
		ram[15'h9DD] =  8'h6E;
		ram[15'h9DE] =  8'h63;
		ram[15'h9DF] =  8'h2C;
		ram[15'h9E0] =  8'h64;
		ram[15'h9E1] =  8'h65;
		ram[15'h9E2] =  8'h63;
		ram[15'h9E3] =  8'h3E;
		ram[15'h9E4] =  8'h20;
		ram[15'h9E5] =  8'h69;
		ram[15'h9E6] =  8'h79;
		ram[15'h9E7] =  8'h2E;
		ram[15'h9E8] =  8'h2E;
		ram[15'h9E9] =  8'h2E;
		ram[15'h9EA] =  8'h2E;
		ram[15'h9EB] =  8'h2E;
		ram[15'h9EC] =  8'h2E;
		ram[15'h9ED] =  8'h2E;
		ram[15'h9EE] =  8'h2E;
		ram[15'h9EF] =  8'h2E;
		ram[15'h9F0] =  8'h2E;
		ram[15'h9F1] =  8'h2E;
		ram[15'h9F2] =  8'h2E;
		ram[15'h9F3] =  8'h2E;
		ram[15'h9F4] =  8'h2E;
		ram[15'h9F5] =  8'h2E;
		ram[15'h9F6] =  8'h2E;
		ram[15'h9F7] =  8'h2E;
		ram[15'h9F8] =  8'h2E;
		ram[15'h9F9] =  8'h24;
		ram[15'h9FA] =  8'hD7;
		ram[15'h9FB] =  8'h2C;
		ram[15'h9FC] =  8'h00;
		ram[15'h9FD] =  8'h00;
		ram[15'h9FE] =  8'h00;
		ram[15'h9FF] =  8'h31;
		ram[15'hA00] =  8'h80;
		ram[15'hA01] =  8'h20;
		ram[15'hA02] =  8'hA5;
		ram[15'hA03] =  8'h56;
		ram[15'hA04] =  8'h43;
		ram[15'hA05] =  8'h09;
		ram[15'hA06] =  8'hB4;
		ram[15'hA07] =  8'hC1;
		ram[15'hA08] =  8'hF4;
		ram[15'hA09] =  8'hA2;
		ram[15'hA0A] =  8'hDF;
		ram[15'hA0B] =  8'hD1;
		ram[15'hA0C] =  8'h3C;
		ram[15'hA0D] =  8'hA2;
		ram[15'hA0E] =  8'h3E;
		ram[15'hA0F] =  8'h01;
		ram[15'hA10] =  8'h00;
		ram[15'hA11] =  8'h00;
		ram[15'hA12] =  8'h00;
		ram[15'hA13] =  8'h00;
		ram[15'hA14] =  8'h00;
		ram[15'hA15] =  8'h00;
		ram[15'hA16] =  8'h00;
		ram[15'hA17] =  8'h00;
		ram[15'hA18] =  8'h00;
		ram[15'hA19] =  8'hFF;
		ram[15'hA1A] =  8'h00;
		ram[15'hA1B] =  8'h00;
		ram[15'hA1C] =  8'h00;
		ram[15'hA1D] =  8'h00;
		ram[15'hA1E] =  8'h00;
		ram[15'hA1F] =  8'h00;
		ram[15'hA20] =  8'h00;
		ram[15'hA21] =  8'h00;
		ram[15'hA22] =  8'h00;
		ram[15'hA23] =  8'h00;
		ram[15'hA24] =  8'h00;
		ram[15'hA25] =  8'h00;
		ram[15'hA26] =  8'h00;
		ram[15'hA27] =  8'h00;
		ram[15'hA28] =  8'h00;
		ram[15'hA29] =  8'h00;
		ram[15'hA2A] =  8'h00;
		ram[15'hA2B] =  8'h00;
		ram[15'hA2C] =  8'h00;
		ram[15'hA2D] =  8'h00;
		ram[15'hA2E] =  8'h00;
		ram[15'hA2F] =  8'h00;
		ram[15'hA30] =  8'h00;
		ram[15'hA31] =  8'h00;
		ram[15'hA32] =  8'h00;
		ram[15'hA33] =  8'hD7;
		ram[15'hA34] =  8'h00;
		ram[15'hA35] =  8'h00;
		ram[15'hA36] =  8'h00;
		ram[15'hA37] =  8'h56;
		ram[15'hA38] =  8'hCD;
		ram[15'hA39] =  8'h06;
		ram[15'hA3A] =  8'hF3;
		ram[15'hA3B] =  8'h3C;
		ram[15'hA3C] =  8'h69;
		ram[15'hA3D] =  8'h6E;
		ram[15'hA3E] =  8'h63;
		ram[15'hA3F] =  8'h2C;
		ram[15'hA40] =  8'h64;
		ram[15'hA41] =  8'h65;
		ram[15'hA42] =  8'h63;
		ram[15'hA43] =  8'h3E;
		ram[15'hA44] =  8'h20;
		ram[15'hA45] =  8'h6C;
		ram[15'hA46] =  8'h2E;
		ram[15'hA47] =  8'h2E;
		ram[15'hA48] =  8'h2E;
		ram[15'hA49] =  8'h2E;
		ram[15'hA4A] =  8'h2E;
		ram[15'hA4B] =  8'h2E;
		ram[15'hA4C] =  8'h2E;
		ram[15'hA4D] =  8'h2E;
		ram[15'hA4E] =  8'h2E;
		ram[15'hA4F] =  8'h2E;
		ram[15'hA50] =  8'h2E;
		ram[15'hA51] =  8'h2E;
		ram[15'hA52] =  8'h2E;
		ram[15'hA53] =  8'h2E;
		ram[15'hA54] =  8'h2E;
		ram[15'hA55] =  8'h2E;
		ram[15'hA56] =  8'h2E;
		ram[15'hA57] =  8'h2E;
		ram[15'hA58] =  8'h2E;
		ram[15'hA59] =  8'h24;
		ram[15'hA5A] =  8'hD7;
		ram[15'hA5B] =  8'h34;
		ram[15'hA5C] =  8'h00;
		ram[15'hA5D] =  8'h00;
		ram[15'hA5E] =  8'h00;
		ram[15'hA5F] =  8'h56;
		ram[15'hA60] =  8'hB8;
		ram[15'hA61] =  8'h7C;
		ram[15'hA62] =  8'h0C;
		ram[15'hA63] =  8'h3E;
		ram[15'hA64] =  8'hE5;
		ram[15'hA65] =  8'h3A;
		ram[15'hA66] =  8'h00;
		ram[15'hA67] =  8'h7E;
		ram[15'hA68] =  8'h87;
		ram[15'hA69] =  8'h58;
		ram[15'hA6A] =  8'hDA;
		ram[15'hA6B] =  8'h15;
		ram[15'hA6C] =  8'h5C;
		ram[15'hA6D] =  8'h37;
		ram[15'hA6E] =  8'h1F;
		ram[15'hA6F] =  8'h01;
		ram[15'hA70] =  8'h00;
		ram[15'hA71] =  8'h00;
		ram[15'hA72] =  8'h00;
		ram[15'hA73] =  8'hFF;
		ram[15'hA74] =  8'h00;
		ram[15'hA75] =  8'h00;
		ram[15'hA76] =  8'h00;
		ram[15'hA77] =  8'h00;
		ram[15'hA78] =  8'h00;
		ram[15'hA79] =  8'h00;
		ram[15'hA7A] =  8'h00;
		ram[15'hA7B] =  8'h00;
		ram[15'hA7C] =  8'h00;
		ram[15'hA7D] =  8'h00;
		ram[15'hA7E] =  8'h00;
		ram[15'hA7F] =  8'h00;
		ram[15'hA80] =  8'h00;
		ram[15'hA81] =  8'h00;
		ram[15'hA82] =  8'h00;
		ram[15'hA83] =  8'h00;
		ram[15'hA84] =  8'h00;
		ram[15'hA85] =  8'h00;
		ram[15'hA86] =  8'h00;
		ram[15'hA87] =  8'h00;
		ram[15'hA88] =  8'h00;
		ram[15'hA89] =  8'h00;
		ram[15'hA8A] =  8'h00;
		ram[15'hA8B] =  8'h00;
		ram[15'hA8C] =  8'h00;
		ram[15'hA8D] =  8'h00;
		ram[15'hA8E] =  8'h00;
		ram[15'hA8F] =  8'h00;
		ram[15'hA90] =  8'h00;
		ram[15'hA91] =  8'h00;
		ram[15'hA92] =  8'h00;
		ram[15'hA93] =  8'hD7;
		ram[15'hA94] =  8'h00;
		ram[15'hA95] =  8'h00;
		ram[15'hA96] =  8'h00;
		ram[15'hA97] =  8'hB8;
		ram[15'hA98] =  8'h3A;
		ram[15'hA99] =  8'hDC;
		ram[15'hA9A] =  8'hEF;
		ram[15'hA9B] =  8'h3C;
		ram[15'hA9C] =  8'h69;
		ram[15'hA9D] =  8'h6E;
		ram[15'hA9E] =  8'h63;
		ram[15'hA9F] =  8'h2C;
		ram[15'hAA0] =  8'h64;
		ram[15'hAA1] =  8'h65;
		ram[15'hAA2] =  8'h63;
		ram[15'hAA3] =  8'h3E;
		ram[15'hAA4] =  8'h20;
		ram[15'hAA5] =  8'h28;
		ram[15'hAA6] =  8'h68;
		ram[15'hAA7] =  8'h6C;
		ram[15'hAA8] =  8'h29;
		ram[15'hAA9] =  8'h2E;
		ram[15'hAAA] =  8'h2E;
		ram[15'hAAB] =  8'h2E;
		ram[15'hAAC] =  8'h2E;
		ram[15'hAAD] =  8'h2E;
		ram[15'hAAE] =  8'h2E;
		ram[15'hAAF] =  8'h2E;
		ram[15'hAB0] =  8'h2E;
		ram[15'hAB1] =  8'h2E;
		ram[15'hAB2] =  8'h2E;
		ram[15'hAB3] =  8'h2E;
		ram[15'hAB4] =  8'h2E;
		ram[15'hAB5] =  8'h2E;
		ram[15'hAB6] =  8'h2E;
		ram[15'hAB7] =  8'h2E;
		ram[15'hAB8] =  8'h2E;
		ram[15'hAB9] =  8'h24;
		ram[15'hABA] =  8'hD7;
		ram[15'hABB] =  8'h33;
		ram[15'hABC] =  8'h00;
		ram[15'hABD] =  8'h00;
		ram[15'hABE] =  8'h00;
		ram[15'hABF] =  8'h6F;
		ram[15'hAC0] =  8'h34;
		ram[15'hAC1] =  8'h82;
		ram[15'hAC2] =  8'hD4;
		ram[15'hAC3] =  8'h69;
		ram[15'hAC4] =  8'hD1;
		ram[15'hAC5] =  8'hB6;
		ram[15'hAC6] =  8'hDE;
		ram[15'hAC7] =  8'h94;
		ram[15'hAC8] =  8'hA4;
		ram[15'hAC9] =  8'h76;
		ram[15'hACA] =  8'hF4;
		ram[15'hACB] =  8'h53;
		ram[15'hACC] =  8'h02;
		ram[15'hACD] =  8'h5B;
		ram[15'hACE] =  8'h85;
		ram[15'hACF] =  8'h08;
		ram[15'hAD0] =  8'h00;
		ram[15'hAD1] =  8'h00;
		ram[15'hAD2] =  8'h00;
		ram[15'hAD3] =  8'h00;
		ram[15'hAD4] =  8'h00;
		ram[15'hAD5] =  8'h00;
		ram[15'hAD6] =  8'h00;
		ram[15'hAD7] =  8'h00;
		ram[15'hAD8] =  8'h00;
		ram[15'hAD9] =  8'h00;
		ram[15'hADA] =  8'h00;
		ram[15'hADB] =  8'h00;
		ram[15'hADC] =  8'h00;
		ram[15'hADD] =  8'h00;
		ram[15'hADE] =  8'h00;
		ram[15'hADF] =  8'h00;
		ram[15'hAE0] =  8'h00;
		ram[15'hAE1] =  8'h21;
		ram[15'hAE2] =  8'hF8;
		ram[15'hAE3] =  8'h00;
		ram[15'hAE4] =  8'h00;
		ram[15'hAE5] =  8'h00;
		ram[15'hAE6] =  8'h00;
		ram[15'hAE7] =  8'h00;
		ram[15'hAE8] =  8'h00;
		ram[15'hAE9] =  8'h00;
		ram[15'hAEA] =  8'h00;
		ram[15'hAEB] =  8'h00;
		ram[15'hAEC] =  8'h00;
		ram[15'hAED] =  8'h00;
		ram[15'hAEE] =  8'h00;
		ram[15'hAEF] =  8'h00;
		ram[15'hAF0] =  8'h00;
		ram[15'hAF1] =  8'h00;
		ram[15'hAF2] =  8'h00;
		ram[15'hAF3] =  8'hD7;
		ram[15'hAF4] =  8'h00;
		ram[15'hAF5] =  8'h00;
		ram[15'hAF6] =  8'h00;
		ram[15'hAF7] =  8'h5D;
		ram[15'hAF8] =  8'hAC;
		ram[15'hAF9] =  8'hD5;
		ram[15'hAFA] =  8'h27;
		ram[15'hAFB] =  8'h3C;
		ram[15'hAFC] =  8'h69;
		ram[15'hAFD] =  8'h6E;
		ram[15'hAFE] =  8'h63;
		ram[15'hAFF] =  8'h2C;
		ram[15'hB00] =  8'h64;
		ram[15'hB01] =  8'h65;
		ram[15'hB02] =  8'h63;
		ram[15'hB03] =  8'h3E;
		ram[15'hB04] =  8'h20;
		ram[15'hB05] =  8'h73;
		ram[15'hB06] =  8'h70;
		ram[15'hB07] =  8'h2E;
		ram[15'hB08] =  8'h2E;
		ram[15'hB09] =  8'h2E;
		ram[15'hB0A] =  8'h2E;
		ram[15'hB0B] =  8'h2E;
		ram[15'hB0C] =  8'h2E;
		ram[15'hB0D] =  8'h2E;
		ram[15'hB0E] =  8'h2E;
		ram[15'hB0F] =  8'h2E;
		ram[15'hB10] =  8'h2E;
		ram[15'hB11] =  8'h2E;
		ram[15'hB12] =  8'h2E;
		ram[15'hB13] =  8'h2E;
		ram[15'hB14] =  8'h2E;
		ram[15'hB15] =  8'h2E;
		ram[15'hB16] =  8'h2E;
		ram[15'hB17] =  8'h2E;
		ram[15'hB18] =  8'h2E;
		ram[15'hB19] =  8'h24;
		ram[15'hB1A] =  8'hD7;
		ram[15'hB1B] =  8'hDD;
		ram[15'hB1C] =  8'h34;
		ram[15'hB1D] =  8'h01;
		ram[15'hB1E] =  8'h00;
		ram[15'hB1F] =  8'h6E;
		ram[15'hB20] =  8'hFA;
		ram[15'hB21] =  8'h39;
		ram[15'hB22] =  8'h00;
		ram[15'hB23] =  8'h39;
		ram[15'hB24] =  8'h00;
		ram[15'hB25] =  8'h28;
		ram[15'hB26] =  8'h2C;
		ram[15'hB27] =  8'h94;
		ram[15'hB28] =  8'h88;
		ram[15'hB29] =  8'h57;
		ram[15'hB2A] =  8'h50;
		ram[15'hB2B] =  8'h16;
		ram[15'hB2C] =  8'h33;
		ram[15'hB2D] =  8'h6F;
		ram[15'hB2E] =  8'h28;
		ram[15'hB2F] =  8'h20;
		ram[15'hB30] =  8'h01;
		ram[15'hB31] =  8'h00;
		ram[15'hB32] =  8'h00;
		ram[15'hB33] =  8'hFF;
		ram[15'hB34] =  8'h00;
		ram[15'hB35] =  8'h00;
		ram[15'hB36] =  8'h00;
		ram[15'hB37] =  8'h00;
		ram[15'hB38] =  8'h00;
		ram[15'hB39] =  8'h00;
		ram[15'hB3A] =  8'h00;
		ram[15'hB3B] =  8'h00;
		ram[15'hB3C] =  8'h00;
		ram[15'hB3D] =  8'h00;
		ram[15'hB3E] =  8'h00;
		ram[15'hB3F] =  8'h00;
		ram[15'hB40] =  8'h00;
		ram[15'hB41] =  8'h00;
		ram[15'hB42] =  8'h00;
		ram[15'hB43] =  8'h00;
		ram[15'hB44] =  8'h00;
		ram[15'hB45] =  8'h00;
		ram[15'hB46] =  8'h00;
		ram[15'hB47] =  8'h00;
		ram[15'hB48] =  8'h00;
		ram[15'hB49] =  8'h00;
		ram[15'hB4A] =  8'h00;
		ram[15'hB4B] =  8'h00;
		ram[15'hB4C] =  8'h00;
		ram[15'hB4D] =  8'h00;
		ram[15'hB4E] =  8'h00;
		ram[15'hB4F] =  8'h00;
		ram[15'hB50] =  8'h00;
		ram[15'hB51] =  8'h00;
		ram[15'hB52] =  8'h00;
		ram[15'hB53] =  8'hD7;
		ram[15'hB54] =  8'h00;
		ram[15'hB55] =  8'h00;
		ram[15'hB56] =  8'h00;
		ram[15'hB57] =  8'h20;
		ram[15'hB58] =  8'h58;
		ram[15'hB59] =  8'h14;
		ram[15'hB5A] =  8'h70;
		ram[15'hB5B] =  8'h3C;
		ram[15'hB5C] =  8'h69;
		ram[15'hB5D] =  8'h6E;
		ram[15'hB5E] =  8'h63;
		ram[15'hB5F] =  8'h2C;
		ram[15'hB60] =  8'h64;
		ram[15'hB61] =  8'h65;
		ram[15'hB62] =  8'h63;
		ram[15'hB63] =  8'h3E;
		ram[15'hB64] =  8'h20;
		ram[15'hB65] =  8'h28;
		ram[15'hB66] =  8'h3C;
		ram[15'hB67] =  8'h69;
		ram[15'hB68] =  8'h78;
		ram[15'hB69] =  8'h2C;
		ram[15'hB6A] =  8'h69;
		ram[15'hB6B] =  8'h79;
		ram[15'hB6C] =  8'h3E;
		ram[15'hB6D] =  8'h2B;
		ram[15'hB6E] =  8'h31;
		ram[15'hB6F] =  8'h29;
		ram[15'hB70] =  8'h2E;
		ram[15'hB71] =  8'h2E;
		ram[15'hB72] =  8'h2E;
		ram[15'hB73] =  8'h2E;
		ram[15'hB74] =  8'h2E;
		ram[15'hB75] =  8'h2E;
		ram[15'hB76] =  8'h2E;
		ram[15'hB77] =  8'h2E;
		ram[15'hB78] =  8'h2E;
		ram[15'hB79] =  8'h24;
		ram[15'hB7A] =  8'hD7;
		ram[15'hB7B] =  8'hDD;
		ram[15'hB7C] =  8'h24;
		ram[15'hB7D] =  8'h00;
		ram[15'hB7E] =  8'h00;
		ram[15'hB7F] =  8'h38;
		ram[15'hB80] =  8'hB8;
		ram[15'hB81] =  8'h6C;
		ram[15'hB82] =  8'h31;
		ram[15'hB83] =  8'hD4;
		ram[15'hB84] =  8'hC6;
		ram[15'hB85] =  8'h01;
		ram[15'hB86] =  8'h3E;
		ram[15'hB87] =  8'h58;
		ram[15'hB88] =  8'h83;
		ram[15'hB89] =  8'hB4;
		ram[15'hB8A] =  8'h15;
		ram[15'hB8B] =  8'h81;
		ram[15'hB8C] =  8'hDE;
		ram[15'hB8D] =  8'h59;
		ram[15'hB8E] =  8'h42;
		ram[15'hB8F] =  8'h00;
		ram[15'hB90] =  8'h01;
		ram[15'hB91] =  8'h00;
		ram[15'hB92] =  8'h00;
		ram[15'hB93] =  8'h00;
		ram[15'hB94] =  8'h00;
		ram[15'hB95] =  8'h00;
		ram[15'hB96] =  8'hFF;
		ram[15'hB97] =  8'h00;
		ram[15'hB98] =  8'h00;
		ram[15'hB99] =  8'h00;
		ram[15'hB9A] =  8'h00;
		ram[15'hB9B] =  8'h00;
		ram[15'hB9C] =  8'h00;
		ram[15'hB9D] =  8'h00;
		ram[15'hB9E] =  8'h00;
		ram[15'hB9F] =  8'h00;
		ram[15'hBA0] =  8'h00;
		ram[15'hBA1] =  8'h00;
		ram[15'hBA2] =  8'h00;
		ram[15'hBA3] =  8'h00;
		ram[15'hBA4] =  8'h00;
		ram[15'hBA5] =  8'h00;
		ram[15'hBA6] =  8'h00;
		ram[15'hBA7] =  8'h00;
		ram[15'hBA8] =  8'h00;
		ram[15'hBA9] =  8'h00;
		ram[15'hBAA] =  8'h00;
		ram[15'hBAB] =  8'h00;
		ram[15'hBAC] =  8'h00;
		ram[15'hBAD] =  8'h00;
		ram[15'hBAE] =  8'h00;
		ram[15'hBAF] =  8'h00;
		ram[15'hBB0] =  8'h00;
		ram[15'hBB1] =  8'h00;
		ram[15'hBB2] =  8'h00;
		ram[15'hBB3] =  8'hD7;
		ram[15'hBB4] =  8'h00;
		ram[15'hBB5] =  8'h00;
		ram[15'hBB6] =  8'h00;
		ram[15'hBB7] =  8'h6F;
		ram[15'hBB8] =  8'h46;
		ram[15'hBB9] =  8'h36;
		ram[15'hBBA] =  8'h62;
		ram[15'hBBB] =  8'h3C;
		ram[15'hBBC] =  8'h69;
		ram[15'hBBD] =  8'h6E;
		ram[15'hBBE] =  8'h63;
		ram[15'hBBF] =  8'h2C;
		ram[15'hBC0] =  8'h64;
		ram[15'hBC1] =  8'h65;
		ram[15'hBC2] =  8'h63;
		ram[15'hBC3] =  8'h3E;
		ram[15'hBC4] =  8'h20;
		ram[15'hBC5] =  8'h69;
		ram[15'hBC6] =  8'h78;
		ram[15'hBC7] =  8'h68;
		ram[15'hBC8] =  8'h2E;
		ram[15'hBC9] =  8'h2E;
		ram[15'hBCA] =  8'h2E;
		ram[15'hBCB] =  8'h2E;
		ram[15'hBCC] =  8'h2E;
		ram[15'hBCD] =  8'h2E;
		ram[15'hBCE] =  8'h2E;
		ram[15'hBCF] =  8'h2E;
		ram[15'hBD0] =  8'h2E;
		ram[15'hBD1] =  8'h2E;
		ram[15'hBD2] =  8'h2E;
		ram[15'hBD3] =  8'h2E;
		ram[15'hBD4] =  8'h2E;
		ram[15'hBD5] =  8'h2E;
		ram[15'hBD6] =  8'h2E;
		ram[15'hBD7] =  8'h2E;
		ram[15'hBD8] =  8'h2E;
		ram[15'hBD9] =  8'h24;
		ram[15'hBDA] =  8'hD7;
		ram[15'hBDB] =  8'hDD;
		ram[15'hBDC] =  8'h2C;
		ram[15'hBDD] =  8'h00;
		ram[15'hBDE] =  8'h00;
		ram[15'hBDF] =  8'h14;
		ram[15'hBE0] =  8'h4D;
		ram[15'hBE1] =  8'h60;
		ram[15'hBE2] =  8'h74;
		ram[15'hBE3] =  8'hD4;
		ram[15'hBE4] =  8'h76;
		ram[15'hBE5] =  8'hE7;
		ram[15'hBE6] =  8'h06;
		ram[15'hBE7] =  8'hA2;
		ram[15'hBE8] =  8'h32;
		ram[15'hBE9] =  8'h3C;
		ram[15'hBEA] =  8'h21;
		ram[15'hBEB] =  8'hD6;
		ram[15'hBEC] =  8'hD7;
		ram[15'hBED] =  8'hA5;
		ram[15'hBEE] =  8'h99;
		ram[15'hBEF] =  8'h00;
		ram[15'hBF0] =  8'h01;
		ram[15'hBF1] =  8'h00;
		ram[15'hBF2] =  8'h00;
		ram[15'hBF3] =  8'h00;
		ram[15'hBF4] =  8'h00;
		ram[15'hBF5] =  8'hFF;
		ram[15'hBF6] =  8'h00;
		ram[15'hBF7] =  8'h00;
		ram[15'hBF8] =  8'h00;
		ram[15'hBF9] =  8'h00;
		ram[15'hBFA] =  8'h00;
		ram[15'hBFB] =  8'h00;
		ram[15'hBFC] =  8'h00;
		ram[15'hBFD] =  8'h00;
		ram[15'hBFE] =  8'h00;
		ram[15'hBFF] =  8'h00;
		ram[15'hC00] =  8'h00;
		ram[15'hC01] =  8'h00;
		ram[15'hC02] =  8'h00;
		ram[15'hC03] =  8'h00;
		ram[15'hC04] =  8'h00;
		ram[15'hC05] =  8'h00;
		ram[15'hC06] =  8'h00;
		ram[15'hC07] =  8'h00;
		ram[15'hC08] =  8'h00;
		ram[15'hC09] =  8'h00;
		ram[15'hC0A] =  8'h00;
		ram[15'hC0B] =  8'h00;
		ram[15'hC0C] =  8'h00;
		ram[15'hC0D] =  8'h00;
		ram[15'hC0E] =  8'h00;
		ram[15'hC0F] =  8'h00;
		ram[15'hC10] =  8'h00;
		ram[15'hC11] =  8'h00;
		ram[15'hC12] =  8'h00;
		ram[15'hC13] =  8'hD7;
		ram[15'hC14] =  8'h00;
		ram[15'hC15] =  8'h00;
		ram[15'hC16] =  8'h00;
		ram[15'hC17] =  8'h02;
		ram[15'hC18] =  8'h7B;
		ram[15'hC19] =  8'hEF;
		ram[15'hC1A] =  8'h2C;
		ram[15'hC1B] =  8'h3C;
		ram[15'hC1C] =  8'h69;
		ram[15'hC1D] =  8'h6E;
		ram[15'hC1E] =  8'h63;
		ram[15'hC1F] =  8'h2C;
		ram[15'hC20] =  8'h64;
		ram[15'hC21] =  8'h65;
		ram[15'hC22] =  8'h63;
		ram[15'hC23] =  8'h3E;
		ram[15'hC24] =  8'h20;
		ram[15'hC25] =  8'h69;
		ram[15'hC26] =  8'h78;
		ram[15'hC27] =  8'h6C;
		ram[15'hC28] =  8'h2E;
		ram[15'hC29] =  8'h2E;
		ram[15'hC2A] =  8'h2E;
		ram[15'hC2B] =  8'h2E;
		ram[15'hC2C] =  8'h2E;
		ram[15'hC2D] =  8'h2E;
		ram[15'hC2E] =  8'h2E;
		ram[15'hC2F] =  8'h2E;
		ram[15'hC30] =  8'h2E;
		ram[15'hC31] =  8'h2E;
		ram[15'hC32] =  8'h2E;
		ram[15'hC33] =  8'h2E;
		ram[15'hC34] =  8'h2E;
		ram[15'hC35] =  8'h2E;
		ram[15'hC36] =  8'h2E;
		ram[15'hC37] =  8'h2E;
		ram[15'hC38] =  8'h2E;
		ram[15'hC39] =  8'h24;
		ram[15'hC3A] =  8'hD7;
		ram[15'hC3B] =  8'hDD;
		ram[15'hC3C] =  8'h24;
		ram[15'hC3D] =  8'h00;
		ram[15'hC3E] =  8'h00;
		ram[15'hC3F] =  8'h36;
		ram[15'hC40] =  8'h28;
		ram[15'hC41] =  8'h6F;
		ram[15'hC42] =  8'h9F;
		ram[15'hC43] =  8'h16;
		ram[15'hC44] =  8'h91;
		ram[15'hC45] =  8'hB9;
		ram[15'hC46] =  8'h61;
		ram[15'hC47] =  8'hCB;
		ram[15'hC48] =  8'h82;
		ram[15'hC49] =  8'h19;
		ram[15'hC4A] =  8'hE2;
		ram[15'hC4B] =  8'h92;
		ram[15'hC4C] =  8'h73;
		ram[15'hC4D] =  8'h8C;
		ram[15'hC4E] =  8'hA9;
		ram[15'hC4F] =  8'h00;
		ram[15'hC50] =  8'h01;
		ram[15'hC51] =  8'h00;
		ram[15'hC52] =  8'h00;
		ram[15'hC53] =  8'h00;
		ram[15'hC54] =  8'hFF;
		ram[15'hC55] =  8'h00;
		ram[15'hC56] =  8'h00;
		ram[15'hC57] =  8'h00;
		ram[15'hC58] =  8'h00;
		ram[15'hC59] =  8'h00;
		ram[15'hC5A] =  8'h00;
		ram[15'hC5B] =  8'h00;
		ram[15'hC5C] =  8'h00;
		ram[15'hC5D] =  8'h00;
		ram[15'hC5E] =  8'h00;
		ram[15'hC5F] =  8'h00;
		ram[15'hC60] =  8'h00;
		ram[15'hC61] =  8'h00;
		ram[15'hC62] =  8'h00;
		ram[15'hC63] =  8'h00;
		ram[15'hC64] =  8'h00;
		ram[15'hC65] =  8'h00;
		ram[15'hC66] =  8'h00;
		ram[15'hC67] =  8'h00;
		ram[15'hC68] =  8'h00;
		ram[15'hC69] =  8'h00;
		ram[15'hC6A] =  8'h00;
		ram[15'hC6B] =  8'h00;
		ram[15'hC6C] =  8'h00;
		ram[15'hC6D] =  8'h00;
		ram[15'hC6E] =  8'h00;
		ram[15'hC6F] =  8'h00;
		ram[15'hC70] =  8'h00;
		ram[15'hC71] =  8'h00;
		ram[15'hC72] =  8'h00;
		ram[15'hC73] =  8'hD7;
		ram[15'hC74] =  8'h00;
		ram[15'hC75] =  8'h00;
		ram[15'hC76] =  8'h00;
		ram[15'hC77] =  8'h2D;
		ram[15'hC78] =  8'h96;
		ram[15'hC79] =  8'h6C;
		ram[15'hC7A] =  8'hF3;
		ram[15'hC7B] =  8'h3C;
		ram[15'hC7C] =  8'h69;
		ram[15'hC7D] =  8'h6E;
		ram[15'hC7E] =  8'h63;
		ram[15'hC7F] =  8'h2C;
		ram[15'hC80] =  8'h64;
		ram[15'hC81] =  8'h65;
		ram[15'hC82] =  8'h63;
		ram[15'hC83] =  8'h3E;
		ram[15'hC84] =  8'h20;
		ram[15'hC85] =  8'h69;
		ram[15'hC86] =  8'h79;
		ram[15'hC87] =  8'h68;
		ram[15'hC88] =  8'h2E;
		ram[15'hC89] =  8'h2E;
		ram[15'hC8A] =  8'h2E;
		ram[15'hC8B] =  8'h2E;
		ram[15'hC8C] =  8'h2E;
		ram[15'hC8D] =  8'h2E;
		ram[15'hC8E] =  8'h2E;
		ram[15'hC8F] =  8'h2E;
		ram[15'hC90] =  8'h2E;
		ram[15'hC91] =  8'h2E;
		ram[15'hC92] =  8'h2E;
		ram[15'hC93] =  8'h2E;
		ram[15'hC94] =  8'h2E;
		ram[15'hC95] =  8'h2E;
		ram[15'hC96] =  8'h2E;
		ram[15'hC97] =  8'h2E;
		ram[15'hC98] =  8'h2E;
		ram[15'hC99] =  8'h24;
		ram[15'hC9A] =  8'hD7;
		ram[15'hC9B] =  8'hDD;
		ram[15'hC9C] =  8'h2C;
		ram[15'hC9D] =  8'h00;
		ram[15'hC9E] =  8'h00;
		ram[15'hC9F] =  8'hC6;
		ram[15'hCA0] =  8'hD7;
		ram[15'hCA1] =  8'hD5;
		ram[15'hCA2] =  8'h62;
		ram[15'hCA3] =  8'h9E;
		ram[15'hCA4] =  8'hA0;
		ram[15'hCA5] =  8'h39;
		ram[15'hCA6] =  8'h70;
		ram[15'hCA7] =  8'h7E;
		ram[15'hCA8] =  8'h3E;
		ram[15'hCA9] =  8'h12;
		ram[15'hCAA] =  8'h9F;
		ram[15'hCAB] =  8'h90;
		ram[15'hCAC] =  8'hD9;
		ram[15'hCAD] =  8'h0F;
		ram[15'hCAE] =  8'h22;
		ram[15'hCAF] =  8'h00;
		ram[15'hCB0] =  8'h01;
		ram[15'hCB1] =  8'h00;
		ram[15'hCB2] =  8'h00;
		ram[15'hCB3] =  8'hFF;
		ram[15'hCB4] =  8'h00;
		ram[15'hCB5] =  8'h00;
		ram[15'hCB6] =  8'h00;
		ram[15'hCB7] =  8'h00;
		ram[15'hCB8] =  8'h00;
		ram[15'hCB9] =  8'h00;
		ram[15'hCBA] =  8'h00;
		ram[15'hCBB] =  8'h00;
		ram[15'hCBC] =  8'h00;
		ram[15'hCBD] =  8'h00;
		ram[15'hCBE] =  8'h00;
		ram[15'hCBF] =  8'h00;
		ram[15'hCC0] =  8'h00;
		ram[15'hCC1] =  8'h00;
		ram[15'hCC2] =  8'h00;
		ram[15'hCC3] =  8'h00;
		ram[15'hCC4] =  8'h00;
		ram[15'hCC5] =  8'h00;
		ram[15'hCC6] =  8'h00;
		ram[15'hCC7] =  8'h00;
		ram[15'hCC8] =  8'h00;
		ram[15'hCC9] =  8'h00;
		ram[15'hCCA] =  8'h00;
		ram[15'hCCB] =  8'h00;
		ram[15'hCCC] =  8'h00;
		ram[15'hCCD] =  8'h00;
		ram[15'hCCE] =  8'h00;
		ram[15'hCCF] =  8'h00;
		ram[15'hCD0] =  8'h00;
		ram[15'hCD1] =  8'h00;
		ram[15'hCD2] =  8'h00;
		ram[15'hCD3] =  8'hD7;
		ram[15'hCD4] =  8'h00;
		ram[15'hCD5] =  8'h00;
		ram[15'hCD6] =  8'h00;
		ram[15'hCD7] =  8'hFB;
		ram[15'hCD8] =  8'hCB;
		ram[15'hCD9] =  8'hBA;
		ram[15'hCDA] =  8'h95;
		ram[15'hCDB] =  8'h3C;
		ram[15'hCDC] =  8'h69;
		ram[15'hCDD] =  8'h6E;
		ram[15'hCDE] =  8'h63;
		ram[15'hCDF] =  8'h2C;
		ram[15'hCE0] =  8'h64;
		ram[15'hCE1] =  8'h65;
		ram[15'hCE2] =  8'h63;
		ram[15'hCE3] =  8'h3E;
		ram[15'hCE4] =  8'h20;
		ram[15'hCE5] =  8'h69;
		ram[15'hCE6] =  8'h79;
		ram[15'hCE7] =  8'h6C;
		ram[15'hCE8] =  8'h2E;
		ram[15'hCE9] =  8'h2E;
		ram[15'hCEA] =  8'h2E;
		ram[15'hCEB] =  8'h2E;
		ram[15'hCEC] =  8'h2E;
		ram[15'hCED] =  8'h2E;
		ram[15'hCEE] =  8'h2E;
		ram[15'hCEF] =  8'h2E;
		ram[15'hCF0] =  8'h2E;
		ram[15'hCF1] =  8'h2E;
		ram[15'hCF2] =  8'h2E;
		ram[15'hCF3] =  8'h2E;
		ram[15'hCF4] =  8'h2E;
		ram[15'hCF5] =  8'h2E;
		ram[15'hCF6] =  8'h2E;
		ram[15'hCF7] =  8'h2E;
		ram[15'hCF8] =  8'h2E;
		ram[15'hCF9] =  8'h24;
		ram[15'hCFA] =  8'hD7;
		ram[15'hCFB] =  8'hED;
		ram[15'hCFC] =  8'h4B;
		ram[15'hCFD] =  8'h3A;
		ram[15'hCFE] =  8'h00;
		ram[15'hCFF] =  8'hA8;
		ram[15'hD00] =  8'hF9;
		ram[15'hD01] =  8'h59;
		ram[15'hD02] =  8'hF5;
		ram[15'hD03] =  8'hA4;
		ram[15'hD04] =  8'h93;
		ram[15'hD05] =  8'hED;
		ram[15'hD06] =  8'hF5;
		ram[15'hD07] =  8'h96;
		ram[15'hD08] =  8'h6F;
		ram[15'hD09] =  8'h68;
		ram[15'hD0A] =  8'hD9;
		ram[15'hD0B] =  8'h86;
		ram[15'hD0C] =  8'hE6;
		ram[15'hD0D] =  8'hD8;
		ram[15'hD0E] =  8'h4B;
		ram[15'hD0F] =  8'h00;
		ram[15'hD10] =  8'h10;
		ram[15'hD11] =  8'h00;
		ram[15'hD12] =  8'h00;
		ram[15'hD13] =  8'h00;
		ram[15'hD14] =  8'h00;
		ram[15'hD15] =  8'h00;
		ram[15'hD16] =  8'h00;
		ram[15'hD17] =  8'h00;
		ram[15'hD18] =  8'h00;
		ram[15'hD19] =  8'h00;
		ram[15'hD1A] =  8'h00;
		ram[15'hD1B] =  8'h00;
		ram[15'hD1C] =  8'h00;
		ram[15'hD1D] =  8'h00;
		ram[15'hD1E] =  8'h00;
		ram[15'hD1F] =  8'h00;
		ram[15'hD20] =  8'h00;
		ram[15'hD21] =  8'h00;
		ram[15'hD22] =  8'h00;
		ram[15'hD23] =  8'h00;
		ram[15'hD24] =  8'h00;
		ram[15'hD25] =  8'h00;
		ram[15'hD26] =  8'h00;
		ram[15'hD27] =  8'hFF;
		ram[15'hD28] =  8'hFF;
		ram[15'hD29] =  8'h00;
		ram[15'hD2A] =  8'h00;
		ram[15'hD2B] =  8'h00;
		ram[15'hD2C] =  8'h00;
		ram[15'hD2D] =  8'h00;
		ram[15'hD2E] =  8'h00;
		ram[15'hD2F] =  8'h00;
		ram[15'hD30] =  8'h00;
		ram[15'hD31] =  8'h00;
		ram[15'hD32] =  8'h00;
		ram[15'hD33] =  8'h00;
		ram[15'hD34] =  8'h00;
		ram[15'hD35] =  8'h00;
		ram[15'hD36] =  8'h00;
		ram[15'hD37] =  8'h4D;
		ram[15'hD38] =  8'h45;
		ram[15'hD39] =  8'hA9;
		ram[15'hD3A] =  8'hAC;
		ram[15'hD3B] =  8'h6C;
		ram[15'hD3C] =  8'h64;
		ram[15'hD3D] =  8'h20;
		ram[15'hD3E] =  8'h3C;
		ram[15'hD3F] =  8'h62;
		ram[15'hD40] =  8'h63;
		ram[15'hD41] =  8'h2C;
		ram[15'hD42] =  8'h64;
		ram[15'hD43] =  8'h65;
		ram[15'hD44] =  8'h3E;
		ram[15'hD45] =  8'h2C;
		ram[15'hD46] =  8'h28;
		ram[15'hD47] =  8'h6E;
		ram[15'hD48] =  8'h6E;
		ram[15'hD49] =  8'h6E;
		ram[15'hD4A] =  8'h6E;
		ram[15'hD4B] =  8'h29;
		ram[15'hD4C] =  8'h2E;
		ram[15'hD4D] =  8'h2E;
		ram[15'hD4E] =  8'h2E;
		ram[15'hD4F] =  8'h2E;
		ram[15'hD50] =  8'h2E;
		ram[15'hD51] =  8'h2E;
		ram[15'hD52] =  8'h2E;
		ram[15'hD53] =  8'h2E;
		ram[15'hD54] =  8'h2E;
		ram[15'hD55] =  8'h2E;
		ram[15'hD56] =  8'h2E;
		ram[15'hD57] =  8'h2E;
		ram[15'hD58] =  8'h2E;
		ram[15'hD59] =  8'h24;
		ram[15'hD5A] =  8'hD7;
		ram[15'hD5B] =  8'h2A;
		ram[15'hD5C] =  8'h3A;
		ram[15'hD5D] =  8'h00;
		ram[15'hD5E] =  8'h00;
		ram[15'hD5F] =  8'h63;
		ram[15'hD60] =  8'h98;
		ram[15'hD61] =  8'h30;
		ram[15'hD62] =  8'h78;
		ram[15'hD63] =  8'h77;
		ram[15'hD64] =  8'h20;
		ram[15'hD65] =  8'hFE;
		ram[15'hD66] =  8'hB1;
		ram[15'hD67] =  8'hFA;
		ram[15'hD68] =  8'hB9;
		ram[15'hD69] =  8'hB8;
		ram[15'hD6A] =  8'hAB;
		ram[15'hD6B] =  8'h04;
		ram[15'hD6C] =  8'h06;
		ram[15'hD6D] =  8'h15;
		ram[15'hD6E] =  8'h60;
		ram[15'hD6F] =  8'h00;
		ram[15'hD70] =  8'h00;
		ram[15'hD71] =  8'h00;
		ram[15'hD72] =  8'h00;
		ram[15'hD73] =  8'h00;
		ram[15'hD74] =  8'h00;
		ram[15'hD75] =  8'h00;
		ram[15'hD76] =  8'h00;
		ram[15'hD77] =  8'h00;
		ram[15'hD78] =  8'h00;
		ram[15'hD79] =  8'h00;
		ram[15'hD7A] =  8'h00;
		ram[15'hD7B] =  8'h00;
		ram[15'hD7C] =  8'h00;
		ram[15'hD7D] =  8'h00;
		ram[15'hD7E] =  8'h00;
		ram[15'hD7F] =  8'h00;
		ram[15'hD80] =  8'h00;
		ram[15'hD81] =  8'h00;
		ram[15'hD82] =  8'h00;
		ram[15'hD83] =  8'h00;
		ram[15'hD84] =  8'h00;
		ram[15'hD85] =  8'h00;
		ram[15'hD86] =  8'h00;
		ram[15'hD87] =  8'hFF;
		ram[15'hD88] =  8'hFF;
		ram[15'hD89] =  8'h00;
		ram[15'hD8A] =  8'h00;
		ram[15'hD8B] =  8'h00;
		ram[15'hD8C] =  8'h00;
		ram[15'hD8D] =  8'h00;
		ram[15'hD8E] =  8'h00;
		ram[15'hD8F] =  8'h00;
		ram[15'hD90] =  8'h00;
		ram[15'hD91] =  8'h00;
		ram[15'hD92] =  8'h00;
		ram[15'hD93] =  8'h00;
		ram[15'hD94] =  8'h00;
		ram[15'hD95] =  8'h00;
		ram[15'hD96] =  8'h00;
		ram[15'hD97] =  8'h5F;
		ram[15'hD98] =  8'h97;
		ram[15'hD99] =  8'h24;
		ram[15'hD9A] =  8'h87;
		ram[15'hD9B] =  8'h6C;
		ram[15'hD9C] =  8'h64;
		ram[15'hD9D] =  8'h20;
		ram[15'hD9E] =  8'h68;
		ram[15'hD9F] =  8'h6C;
		ram[15'hDA0] =  8'h2C;
		ram[15'hDA1] =  8'h28;
		ram[15'hDA2] =  8'h6E;
		ram[15'hDA3] =  8'h6E;
		ram[15'hDA4] =  8'h6E;
		ram[15'hDA5] =  8'h6E;
		ram[15'hDA6] =  8'h29;
		ram[15'hDA7] =  8'h2E;
		ram[15'hDA8] =  8'h2E;
		ram[15'hDA9] =  8'h2E;
		ram[15'hDAA] =  8'h2E;
		ram[15'hDAB] =  8'h2E;
		ram[15'hDAC] =  8'h2E;
		ram[15'hDAD] =  8'h2E;
		ram[15'hDAE] =  8'h2E;
		ram[15'hDAF] =  8'h2E;
		ram[15'hDB0] =  8'h2E;
		ram[15'hDB1] =  8'h2E;
		ram[15'hDB2] =  8'h2E;
		ram[15'hDB3] =  8'h2E;
		ram[15'hDB4] =  8'h2E;
		ram[15'hDB5] =  8'h2E;
		ram[15'hDB6] =  8'h2E;
		ram[15'hDB7] =  8'h2E;
		ram[15'hDB8] =  8'h2E;
		ram[15'hDB9] =  8'h24;
		ram[15'hDBA] =  8'hD7;
		ram[15'hDBB] =  8'hED;
		ram[15'hDBC] =  8'h7B;
		ram[15'hDBD] =  8'h3A;
		ram[15'hDBE] =  8'h00;
		ram[15'hDBF] =  8'hFC;
		ram[15'hDC0] =  8'h8D;
		ram[15'hDC1] =  8'hD7;
		ram[15'hDC2] =  8'h57;
		ram[15'hDC3] =  8'h61;
		ram[15'hDC4] =  8'h21;
		ram[15'hDC5] =  8'h18;
		ram[15'hDC6] =  8'hCA;
		ram[15'hDC7] =  8'h85;
		ram[15'hDC8] =  8'hC1;
		ram[15'hDC9] =  8'hDA;
		ram[15'hDCA] =  8'h27;
		ram[15'hDCB] =  8'h83;
		ram[15'hDCC] =  8'h1E;
		ram[15'hDCD] =  8'h60;
		ram[15'hDCE] =  8'hF4;
		ram[15'hDCF] =  8'h00;
		ram[15'hDD0] =  8'h00;
		ram[15'hDD1] =  8'h00;
		ram[15'hDD2] =  8'h00;
		ram[15'hDD3] =  8'h00;
		ram[15'hDD4] =  8'h00;
		ram[15'hDD5] =  8'h00;
		ram[15'hDD6] =  8'h00;
		ram[15'hDD7] =  8'h00;
		ram[15'hDD8] =  8'h00;
		ram[15'hDD9] =  8'h00;
		ram[15'hDDA] =  8'h00;
		ram[15'hDDB] =  8'h00;
		ram[15'hDDC] =  8'h00;
		ram[15'hDDD] =  8'h00;
		ram[15'hDDE] =  8'h00;
		ram[15'hDDF] =  8'h00;
		ram[15'hDE0] =  8'h00;
		ram[15'hDE1] =  8'h00;
		ram[15'hDE2] =  8'h00;
		ram[15'hDE3] =  8'h00;
		ram[15'hDE4] =  8'h00;
		ram[15'hDE5] =  8'h00;
		ram[15'hDE6] =  8'h00;
		ram[15'hDE7] =  8'hFF;
		ram[15'hDE8] =  8'hFF;
		ram[15'hDE9] =  8'h00;
		ram[15'hDEA] =  8'h00;
		ram[15'hDEB] =  8'h00;
		ram[15'hDEC] =  8'h00;
		ram[15'hDED] =  8'h00;
		ram[15'hDEE] =  8'h00;
		ram[15'hDEF] =  8'h00;
		ram[15'hDF0] =  8'h00;
		ram[15'hDF1] =  8'h00;
		ram[15'hDF2] =  8'h00;
		ram[15'hDF3] =  8'h00;
		ram[15'hDF4] =  8'h00;
		ram[15'hDF5] =  8'h00;
		ram[15'hDF6] =  8'h00;
		ram[15'hDF7] =  8'h7A;
		ram[15'hDF8] =  8'hCE;
		ram[15'hDF9] =  8'hA1;
		ram[15'hDFA] =  8'h1B;
		ram[15'hDFB] =  8'h6C;
		ram[15'hDFC] =  8'h64;
		ram[15'hDFD] =  8'h20;
		ram[15'hDFE] =  8'h73;
		ram[15'hDFF] =  8'h70;
		ram[15'hE00] =  8'h2C;
		ram[15'hE01] =  8'h28;
		ram[15'hE02] =  8'h6E;
		ram[15'hE03] =  8'h6E;
		ram[15'hE04] =  8'h6E;
		ram[15'hE05] =  8'h6E;
		ram[15'hE06] =  8'h29;
		ram[15'hE07] =  8'h2E;
		ram[15'hE08] =  8'h2E;
		ram[15'hE09] =  8'h2E;
		ram[15'hE0A] =  8'h2E;
		ram[15'hE0B] =  8'h2E;
		ram[15'hE0C] =  8'h2E;
		ram[15'hE0D] =  8'h2E;
		ram[15'hE0E] =  8'h2E;
		ram[15'hE0F] =  8'h2E;
		ram[15'hE10] =  8'h2E;
		ram[15'hE11] =  8'h2E;
		ram[15'hE12] =  8'h2E;
		ram[15'hE13] =  8'h2E;
		ram[15'hE14] =  8'h2E;
		ram[15'hE15] =  8'h2E;
		ram[15'hE16] =  8'h2E;
		ram[15'hE17] =  8'h2E;
		ram[15'hE18] =  8'h2E;
		ram[15'hE19] =  8'h24;
		ram[15'hE1A] =  8'hD7;
		ram[15'hE1B] =  8'hDD;
		ram[15'hE1C] =  8'h2A;
		ram[15'hE1D] =  8'h3A;
		ram[15'hE1E] =  8'h00;
		ram[15'hE1F] =  8'hD7;
		ram[15'hE20] =  8'hDE;
		ram[15'hE21] =  8'hFA;
		ram[15'hE22] =  8'hA6;
		ram[15'hE23] =  8'h80;
		ram[15'hE24] =  8'hF7;
		ram[15'hE25] =  8'h4C;
		ram[15'hE26] =  8'h24;
		ram[15'hE27] =  8'hDE;
		ram[15'hE28] =  8'h87;
		ram[15'hE29] =  8'hC2;
		ram[15'hE2A] =  8'hBC;
		ram[15'hE2B] =  8'h16;
		ram[15'hE2C] =  8'h63;
		ram[15'hE2D] =  8'h96;
		ram[15'hE2E] =  8'h4C;
		ram[15'hE2F] =  8'h20;
		ram[15'hE30] =  8'h00;
		ram[15'hE31] =  8'h00;
		ram[15'hE32] =  8'h00;
		ram[15'hE33] =  8'h00;
		ram[15'hE34] =  8'h00;
		ram[15'hE35] =  8'h00;
		ram[15'hE36] =  8'h00;
		ram[15'hE37] =  8'h00;
		ram[15'hE38] =  8'h00;
		ram[15'hE39] =  8'h00;
		ram[15'hE3A] =  8'h00;
		ram[15'hE3B] =  8'h00;
		ram[15'hE3C] =  8'h00;
		ram[15'hE3D] =  8'h00;
		ram[15'hE3E] =  8'h00;
		ram[15'hE3F] =  8'h00;
		ram[15'hE40] =  8'h00;
		ram[15'hE41] =  8'h00;
		ram[15'hE42] =  8'h00;
		ram[15'hE43] =  8'h00;
		ram[15'hE44] =  8'h00;
		ram[15'hE45] =  8'h00;
		ram[15'hE46] =  8'h00;
		ram[15'hE47] =  8'hFF;
		ram[15'hE48] =  8'hFF;
		ram[15'hE49] =  8'h00;
		ram[15'hE4A] =  8'h00;
		ram[15'hE4B] =  8'h00;
		ram[15'hE4C] =  8'h00;
		ram[15'hE4D] =  8'h00;
		ram[15'hE4E] =  8'h00;
		ram[15'hE4F] =  8'h00;
		ram[15'hE50] =  8'h00;
		ram[15'hE51] =  8'h00;
		ram[15'hE52] =  8'h00;
		ram[15'hE53] =  8'h00;
		ram[15'hE54] =  8'h00;
		ram[15'hE55] =  8'h00;
		ram[15'hE56] =  8'h00;
		ram[15'hE57] =  8'h85;
		ram[15'hE58] =  8'h8B;
		ram[15'hE59] =  8'hF1;
		ram[15'hE5A] =  8'h6D;
		ram[15'hE5B] =  8'h6C;
		ram[15'hE5C] =  8'h64;
		ram[15'hE5D] =  8'h20;
		ram[15'hE5E] =  8'h3C;
		ram[15'hE5F] =  8'h69;
		ram[15'hE60] =  8'h78;
		ram[15'hE61] =  8'h2C;
		ram[15'hE62] =  8'h69;
		ram[15'hE63] =  8'h79;
		ram[15'hE64] =  8'h3E;
		ram[15'hE65] =  8'h2C;
		ram[15'hE66] =  8'h28;
		ram[15'hE67] =  8'h6E;
		ram[15'hE68] =  8'h6E;
		ram[15'hE69] =  8'h6E;
		ram[15'hE6A] =  8'h6E;
		ram[15'hE6B] =  8'h29;
		ram[15'hE6C] =  8'h2E;
		ram[15'hE6D] =  8'h2E;
		ram[15'hE6E] =  8'h2E;
		ram[15'hE6F] =  8'h2E;
		ram[15'hE70] =  8'h2E;
		ram[15'hE71] =  8'h2E;
		ram[15'hE72] =  8'h2E;
		ram[15'hE73] =  8'h2E;
		ram[15'hE74] =  8'h2E;
		ram[15'hE75] =  8'h2E;
		ram[15'hE76] =  8'h2E;
		ram[15'hE77] =  8'h2E;
		ram[15'hE78] =  8'h2E;
		ram[15'hE79] =  8'h24;
		ram[15'hE7A] =  8'hD7;
		ram[15'hE7B] =  8'hED;
		ram[15'hE7C] =  8'h43;
		ram[15'hE7D] =  8'h3A;
		ram[15'hE7E] =  8'h00;
		ram[15'hE7F] =  8'h98;
		ram[15'hE80] =  8'h1F;
		ram[15'hE81] =  8'h4D;
		ram[15'hE82] =  8'h84;
		ram[15'hE83] =  8'hAC;
		ram[15'hE84] =  8'hE8;
		ram[15'hE85] =  8'hED;
		ram[15'hE86] =  8'hC9;
		ram[15'hE87] =  8'h5D;
		ram[15'hE88] =  8'hC9;
		ram[15'hE89] =  8'h61;
		ram[15'hE8A] =  8'h8F;
		ram[15'hE8B] =  8'h80;
		ram[15'hE8C] =  8'h3F;
		ram[15'hE8D] =  8'hBF;
		ram[15'hE8E] =  8'hC7;
		ram[15'hE8F] =  8'h00;
		ram[15'hE90] =  8'h10;
		ram[15'hE91] =  8'h00;
		ram[15'hE92] =  8'h00;
		ram[15'hE93] =  8'h00;
		ram[15'hE94] =  8'h00;
		ram[15'hE95] =  8'h00;
		ram[15'hE96] =  8'h00;
		ram[15'hE97] =  8'h00;
		ram[15'hE98] =  8'h00;
		ram[15'hE99] =  8'h00;
		ram[15'hE9A] =  8'h00;
		ram[15'hE9B] =  8'h00;
		ram[15'hE9C] =  8'h00;
		ram[15'hE9D] =  8'h00;
		ram[15'hE9E] =  8'h00;
		ram[15'hE9F] =  8'h00;
		ram[15'hEA0] =  8'h00;
		ram[15'hEA1] =  8'h00;
		ram[15'hEA2] =  8'h00;
		ram[15'hEA3] =  8'h00;
		ram[15'hEA4] =  8'h00;
		ram[15'hEA5] =  8'h00;
		ram[15'hEA6] =  8'h00;
		ram[15'hEA7] =  8'h00;
		ram[15'hEA8] =  8'h00;
		ram[15'hEA9] =  8'h00;
		ram[15'hEAA] =  8'h00;
		ram[15'hEAB] =  8'h00;
		ram[15'hEAC] =  8'h00;
		ram[15'hEAD] =  8'h00;
		ram[15'hEAE] =  8'h00;
		ram[15'hEAF] =  8'hFF;
		ram[15'hEB0] =  8'hFF;
		ram[15'hEB1] =  8'hFF;
		ram[15'hEB2] =  8'hFF;
		ram[15'hEB3] =  8'h00;
		ram[15'hEB4] =  8'h00;
		ram[15'hEB5] =  8'h00;
		ram[15'hEB6] =  8'h00;
		ram[15'hEB7] =  8'h64;
		ram[15'hEB8] =  8'h1E;
		ram[15'hEB9] =  8'h87;
		ram[15'hEBA] =  8'h15;
		ram[15'hEBB] =  8'h6C;
		ram[15'hEBC] =  8'h64;
		ram[15'hEBD] =  8'h20;
		ram[15'hEBE] =  8'h28;
		ram[15'hEBF] =  8'h6E;
		ram[15'hEC0] =  8'h6E;
		ram[15'hEC1] =  8'h6E;
		ram[15'hEC2] =  8'h6E;
		ram[15'hEC3] =  8'h29;
		ram[15'hEC4] =  8'h2C;
		ram[15'hEC5] =  8'h3C;
		ram[15'hEC6] =  8'h62;
		ram[15'hEC7] =  8'h63;
		ram[15'hEC8] =  8'h2C;
		ram[15'hEC9] =  8'h64;
		ram[15'hECA] =  8'h65;
		ram[15'hECB] =  8'h3E;
		ram[15'hECC] =  8'h2E;
		ram[15'hECD] =  8'h2E;
		ram[15'hECE] =  8'h2E;
		ram[15'hECF] =  8'h2E;
		ram[15'hED0] =  8'h2E;
		ram[15'hED1] =  8'h2E;
		ram[15'hED2] =  8'h2E;
		ram[15'hED3] =  8'h2E;
		ram[15'hED4] =  8'h2E;
		ram[15'hED5] =  8'h2E;
		ram[15'hED6] =  8'h2E;
		ram[15'hED7] =  8'h2E;
		ram[15'hED8] =  8'h2E;
		ram[15'hED9] =  8'h24;
		ram[15'hEDA] =  8'hD7;
		ram[15'hEDB] =  8'h22;
		ram[15'hEDC] =  8'h3A;
		ram[15'hEDD] =  8'h00;
		ram[15'hEDE] =  8'h00;
		ram[15'hEDF] =  8'h03;
		ram[15'hEE0] =  8'hD0;
		ram[15'hEE1] =  8'h72;
		ram[15'hEE2] =  8'h77;
		ram[15'hEE3] =  8'h53;
		ram[15'hEE4] =  8'h7F;
		ram[15'hEE5] =  8'h72;
		ram[15'hEE6] =  8'h3F;
		ram[15'hEE7] =  8'hEA;
		ram[15'hEE8] =  8'h64;
		ram[15'hEE9] =  8'h80;
		ram[15'hEEA] =  8'hE1;
		ram[15'hEEB] =  8'h10;
		ram[15'hEEC] =  8'h2D;
		ram[15'hEED] =  8'hE9;
		ram[15'hEEE] =  8'h35;
		ram[15'hEEF] =  8'h00;
		ram[15'hEF0] =  8'h00;
		ram[15'hEF1] =  8'h00;
		ram[15'hEF2] =  8'h00;
		ram[15'hEF3] =  8'h00;
		ram[15'hEF4] =  8'h00;
		ram[15'hEF5] =  8'h00;
		ram[15'hEF6] =  8'h00;
		ram[15'hEF7] =  8'h00;
		ram[15'hEF8] =  8'h00;
		ram[15'hEF9] =  8'h00;
		ram[15'hEFA] =  8'h00;
		ram[15'hEFB] =  8'h00;
		ram[15'hEFC] =  8'h00;
		ram[15'hEFD] =  8'h00;
		ram[15'hEFE] =  8'h00;
		ram[15'hEFF] =  8'h00;
		ram[15'hF00] =  8'h00;
		ram[15'hF01] =  8'h00;
		ram[15'hF02] =  8'h00;
		ram[15'hF03] =  8'h00;
		ram[15'hF04] =  8'h00;
		ram[15'hF05] =  8'h00;
		ram[15'hF06] =  8'h00;
		ram[15'hF07] =  8'h00;
		ram[15'hF08] =  8'h00;
		ram[15'hF09] =  8'h00;
		ram[15'hF0A] =  8'h00;
		ram[15'hF0B] =  8'h00;
		ram[15'hF0C] =  8'h00;
		ram[15'hF0D] =  8'hFF;
		ram[15'hF0E] =  8'hFF;
		ram[15'hF0F] =  8'h00;
		ram[15'hF10] =  8'h00;
		ram[15'hF11] =  8'h00;
		ram[15'hF12] =  8'h00;
		ram[15'hF13] =  8'h00;
		ram[15'hF14] =  8'h00;
		ram[15'hF15] =  8'h00;
		ram[15'hF16] =  8'h00;
		ram[15'hF17] =  8'hA3;
		ram[15'hF18] =  8'h60;
		ram[15'hF19] =  8'h8B;
		ram[15'hF1A] =  8'h47;
		ram[15'hF1B] =  8'h6C;
		ram[15'hF1C] =  8'h64;
		ram[15'hF1D] =  8'h20;
		ram[15'hF1E] =  8'h28;
		ram[15'hF1F] =  8'h6E;
		ram[15'hF20] =  8'h6E;
		ram[15'hF21] =  8'h6E;
		ram[15'hF22] =  8'h6E;
		ram[15'hF23] =  8'h29;
		ram[15'hF24] =  8'h2C;
		ram[15'hF25] =  8'h68;
		ram[15'hF26] =  8'h6C;
		ram[15'hF27] =  8'h2E;
		ram[15'hF28] =  8'h2E;
		ram[15'hF29] =  8'h2E;
		ram[15'hF2A] =  8'h2E;
		ram[15'hF2B] =  8'h2E;
		ram[15'hF2C] =  8'h2E;
		ram[15'hF2D] =  8'h2E;
		ram[15'hF2E] =  8'h2E;
		ram[15'hF2F] =  8'h2E;
		ram[15'hF30] =  8'h2E;
		ram[15'hF31] =  8'h2E;
		ram[15'hF32] =  8'h2E;
		ram[15'hF33] =  8'h2E;
		ram[15'hF34] =  8'h2E;
		ram[15'hF35] =  8'h2E;
		ram[15'hF36] =  8'h2E;
		ram[15'hF37] =  8'h2E;
		ram[15'hF38] =  8'h2E;
		ram[15'hF39] =  8'h24;
		ram[15'hF3A] =  8'hD7;
		ram[15'hF3B] =  8'hED;
		ram[15'hF3C] =  8'h73;
		ram[15'hF3D] =  8'h3A;
		ram[15'hF3E] =  8'h00;
		ram[15'hF3F] =  8'hDC;
		ram[15'hF40] =  8'hC0;
		ram[15'hF41] =  8'hD6;
		ram[15'hF42] =  8'hD1;
		ram[15'hF43] =  8'h5A;
		ram[15'hF44] =  8'hED;
		ram[15'hF45] =  8'h56;
		ram[15'hF46] =  8'hF3;
		ram[15'hF47] =  8'hDA;
		ram[15'hF48] =  8'hAF;
		ram[15'hF49] =  8'hA7;
		ram[15'hF4A] =  8'h6C;
		ram[15'hF4B] =  8'h44;
		ram[15'hF4C] =  8'h9F;
		ram[15'hF4D] =  8'h0A;
		ram[15'hF4E] =  8'h3F;
		ram[15'hF4F] =  8'h00;
		ram[15'hF50] =  8'h00;
		ram[15'hF51] =  8'h00;
		ram[15'hF52] =  8'h00;
		ram[15'hF53] =  8'h00;
		ram[15'hF54] =  8'h00;
		ram[15'hF55] =  8'h00;
		ram[15'hF56] =  8'h00;
		ram[15'hF57] =  8'h00;
		ram[15'hF58] =  8'h00;
		ram[15'hF59] =  8'h00;
		ram[15'hF5A] =  8'h00;
		ram[15'hF5B] =  8'h00;
		ram[15'hF5C] =  8'h00;
		ram[15'hF5D] =  8'h00;
		ram[15'hF5E] =  8'h00;
		ram[15'hF5F] =  8'h00;
		ram[15'hF60] =  8'h00;
		ram[15'hF61] =  8'h00;
		ram[15'hF62] =  8'h00;
		ram[15'hF63] =  8'h00;
		ram[15'hF64] =  8'h00;
		ram[15'hF65] =  8'h00;
		ram[15'hF66] =  8'h00;
		ram[15'hF67] =  8'h00;
		ram[15'hF68] =  8'h00;
		ram[15'hF69] =  8'h00;
		ram[15'hF6A] =  8'h00;
		ram[15'hF6B] =  8'h00;
		ram[15'hF6C] =  8'h00;
		ram[15'hF6D] =  8'h00;
		ram[15'hF6E] =  8'h00;
		ram[15'hF6F] =  8'h00;
		ram[15'hF70] =  8'h00;
		ram[15'hF71] =  8'h00;
		ram[15'hF72] =  8'h00;
		ram[15'hF73] =  8'h00;
		ram[15'hF74] =  8'h00;
		ram[15'hF75] =  8'hFF;
		ram[15'hF76] =  8'hFF;
		ram[15'hF77] =  8'h16;
		ram[15'hF78] =  8'h58;
		ram[15'hF79] =  8'h5F;
		ram[15'hF7A] =  8'hD7;
		ram[15'hF7B] =  8'h6C;
		ram[15'hF7C] =  8'h64;
		ram[15'hF7D] =  8'h20;
		ram[15'hF7E] =  8'h28;
		ram[15'hF7F] =  8'h6E;
		ram[15'hF80] =  8'h6E;
		ram[15'hF81] =  8'h6E;
		ram[15'hF82] =  8'h6E;
		ram[15'hF83] =  8'h29;
		ram[15'hF84] =  8'h2C;
		ram[15'hF85] =  8'h73;
		ram[15'hF86] =  8'h70;
		ram[15'hF87] =  8'h2E;
		ram[15'hF88] =  8'h2E;
		ram[15'hF89] =  8'h2E;
		ram[15'hF8A] =  8'h2E;
		ram[15'hF8B] =  8'h2E;
		ram[15'hF8C] =  8'h2E;
		ram[15'hF8D] =  8'h2E;
		ram[15'hF8E] =  8'h2E;
		ram[15'hF8F] =  8'h2E;
		ram[15'hF90] =  8'h2E;
		ram[15'hF91] =  8'h2E;
		ram[15'hF92] =  8'h2E;
		ram[15'hF93] =  8'h2E;
		ram[15'hF94] =  8'h2E;
		ram[15'hF95] =  8'h2E;
		ram[15'hF96] =  8'h2E;
		ram[15'hF97] =  8'h2E;
		ram[15'hF98] =  8'h2E;
		ram[15'hF99] =  8'h24;
		ram[15'hF9A] =  8'hD7;
		ram[15'hF9B] =  8'hDD;
		ram[15'hF9C] =  8'h22;
		ram[15'hF9D] =  8'h3A;
		ram[15'hF9E] =  8'h00;
		ram[15'hF9F] =  8'hC3;
		ram[15'hFA0] =  8'h6C;
		ram[15'hFA1] =  8'h91;
		ram[15'hFA2] =  8'h0D;
		ram[15'hFA3] =  8'h00;
		ram[15'hFA4] =  8'h69;
		ram[15'hFA5] =  8'hF8;
		ram[15'hFA6] =  8'h8E;
		ram[15'hFA7] =  8'hD6;
		ram[15'hFA8] =  8'hE3;
		ram[15'hFA9] =  8'hF7;
		ram[15'hFAA] =  8'hC3;
		ram[15'hFAB] =  8'hC6;
		ram[15'hFAC] =  8'hD9;
		ram[15'hFAD] =  8'hDF;
		ram[15'hFAE] =  8'hC2;
		ram[15'hFAF] =  8'h20;
		ram[15'hFB0] =  8'h00;
		ram[15'hFB1] =  8'h00;
		ram[15'hFB2] =  8'h00;
		ram[15'hFB3] =  8'h00;
		ram[15'hFB4] =  8'h00;
		ram[15'hFB5] =  8'h00;
		ram[15'hFB6] =  8'h00;
		ram[15'hFB7] =  8'h00;
		ram[15'hFB8] =  8'h00;
		ram[15'hFB9] =  8'h00;
		ram[15'hFBA] =  8'h00;
		ram[15'hFBB] =  8'h00;
		ram[15'hFBC] =  8'h00;
		ram[15'hFBD] =  8'h00;
		ram[15'hFBE] =  8'h00;
		ram[15'hFBF] =  8'h00;
		ram[15'hFC0] =  8'h00;
		ram[15'hFC1] =  8'h00;
		ram[15'hFC2] =  8'h00;
		ram[15'hFC3] =  8'h00;
		ram[15'hFC4] =  8'h00;
		ram[15'hFC5] =  8'h00;
		ram[15'hFC6] =  8'h00;
		ram[15'hFC7] =  8'h00;
		ram[15'hFC8] =  8'h00;
		ram[15'hFC9] =  8'hFF;
		ram[15'hFCA] =  8'hFF;
		ram[15'hFCB] =  8'hFF;
		ram[15'hFCC] =  8'hFF;
		ram[15'hFCD] =  8'h00;
		ram[15'hFCE] =  8'h00;
		ram[15'hFCF] =  8'h00;
		ram[15'hFD0] =  8'h00;
		ram[15'hFD1] =  8'h00;
		ram[15'hFD2] =  8'h00;
		ram[15'hFD3] =  8'h00;
		ram[15'hFD4] =  8'h00;
		ram[15'hFD5] =  8'h00;
		ram[15'hFD6] =  8'h00;
		ram[15'hFD7] =  8'hBA;
		ram[15'hFD8] =  8'h10;
		ram[15'hFD9] =  8'h2A;
		ram[15'hFDA] =  8'h6B;
		ram[15'hFDB] =  8'h6C;
		ram[15'hFDC] =  8'h64;
		ram[15'hFDD] =  8'h20;
		ram[15'hFDE] =  8'h28;
		ram[15'hFDF] =  8'h6E;
		ram[15'hFE0] =  8'h6E;
		ram[15'hFE1] =  8'h6E;
		ram[15'hFE2] =  8'h6E;
		ram[15'hFE3] =  8'h29;
		ram[15'hFE4] =  8'h2C;
		ram[15'hFE5] =  8'h3C;
		ram[15'hFE6] =  8'h69;
		ram[15'hFE7] =  8'h78;
		ram[15'hFE8] =  8'h2C;
		ram[15'hFE9] =  8'h69;
		ram[15'hFEA] =  8'h79;
		ram[15'hFEB] =  8'h3E;
		ram[15'hFEC] =  8'h2E;
		ram[15'hFED] =  8'h2E;
		ram[15'hFEE] =  8'h2E;
		ram[15'hFEF] =  8'h2E;
		ram[15'hFF0] =  8'h2E;
		ram[15'hFF1] =  8'h2E;
		ram[15'hFF2] =  8'h2E;
		ram[15'hFF3] =  8'h2E;
		ram[15'hFF4] =  8'h2E;
		ram[15'hFF5] =  8'h2E;
		ram[15'hFF6] =  8'h2E;
		ram[15'hFF7] =  8'h2E;
		ram[15'hFF8] =  8'h2E;
		ram[15'hFF9] =  8'h24;
		ram[15'hFFA] =  8'hD7;
		ram[15'hFFB] =  8'h01;
		ram[15'hFFC] =  8'h00;
		ram[15'hFFD] =  8'h00;
		ram[15'hFFE] =  8'h00;
		ram[15'hFFF] =  8'h1C;
		ram[15'h1000] =  8'h5C;
		ram[15'h1001] =  8'h46;
		ram[15'h1002] =  8'h2D;
		ram[15'h1003] =  8'hB9;
		ram[15'h1004] =  8'h8E;
		ram[15'h1005] =  8'h78;
		ram[15'h1006] =  8'h60;
		ram[15'h1007] =  8'hB1;
		ram[15'h1008] =  8'h74;
		ram[15'h1009] =  8'h0E;
		ram[15'h100A] =  8'hB3;
		ram[15'h100B] =  8'h46;
		ram[15'h100C] =  8'hD1;
		ram[15'h100D] =  8'hCC;
		ram[15'h100E] =  8'h30;
		ram[15'h100F] =  8'h30;
		ram[15'h1010] =  8'h00;
		ram[15'h1011] =  8'h00;
		ram[15'h1012] =  8'h00;
		ram[15'h1013] =  8'h00;
		ram[15'h1014] =  8'h00;
		ram[15'h1015] =  8'h00;
		ram[15'h1016] =  8'h00;
		ram[15'h1017] =  8'h00;
		ram[15'h1018] =  8'h00;
		ram[15'h1019] =  8'h00;
		ram[15'h101A] =  8'h00;
		ram[15'h101B] =  8'h00;
		ram[15'h101C] =  8'h00;
		ram[15'h101D] =  8'h00;
		ram[15'h101E] =  8'h00;
		ram[15'h101F] =  8'h00;
		ram[15'h1020] =  8'h00;
		ram[15'h1021] =  8'h00;
		ram[15'h1022] =  8'h00;
		ram[15'h1023] =  8'h00;
		ram[15'h1024] =  8'hFF;
		ram[15'h1025] =  8'hFF;
		ram[15'h1026] =  8'h00;
		ram[15'h1027] =  8'h00;
		ram[15'h1028] =  8'h00;
		ram[15'h1029] =  8'h00;
		ram[15'h102A] =  8'h00;
		ram[15'h102B] =  8'h00;
		ram[15'h102C] =  8'h00;
		ram[15'h102D] =  8'h00;
		ram[15'h102E] =  8'h00;
		ram[15'h102F] =  8'h00;
		ram[15'h1030] =  8'h00;
		ram[15'h1031] =  8'h00;
		ram[15'h1032] =  8'h00;
		ram[15'h1033] =  8'h00;
		ram[15'h1034] =  8'h00;
		ram[15'h1035] =  8'h00;
		ram[15'h1036] =  8'h00;
		ram[15'h1037] =  8'hDE;
		ram[15'h1038] =  8'h39;
		ram[15'h1039] =  8'h19;
		ram[15'h103A] =  8'h69;
		ram[15'h103B] =  8'h6C;
		ram[15'h103C] =  8'h64;
		ram[15'h103D] =  8'h20;
		ram[15'h103E] =  8'h3C;
		ram[15'h103F] =  8'h62;
		ram[15'h1040] =  8'h63;
		ram[15'h1041] =  8'h2C;
		ram[15'h1042] =  8'h64;
		ram[15'h1043] =  8'h65;
		ram[15'h1044] =  8'h2C;
		ram[15'h1045] =  8'h68;
		ram[15'h1046] =  8'h6C;
		ram[15'h1047] =  8'h2C;
		ram[15'h1048] =  8'h73;
		ram[15'h1049] =  8'h70;
		ram[15'h104A] =  8'h3E;
		ram[15'h104B] =  8'h2C;
		ram[15'h104C] =  8'h6E;
		ram[15'h104D] =  8'h6E;
		ram[15'h104E] =  8'h6E;
		ram[15'h104F] =  8'h6E;
		ram[15'h1050] =  8'h2E;
		ram[15'h1051] =  8'h2E;
		ram[15'h1052] =  8'h2E;
		ram[15'h1053] =  8'h2E;
		ram[15'h1054] =  8'h2E;
		ram[15'h1055] =  8'h2E;
		ram[15'h1056] =  8'h2E;
		ram[15'h1057] =  8'h2E;
		ram[15'h1058] =  8'h2E;
		ram[15'h1059] =  8'h24;
		ram[15'h105A] =  8'hD7;
		ram[15'h105B] =  8'hDD;
		ram[15'h105C] =  8'h21;
		ram[15'h105D] =  8'h00;
		ram[15'h105E] =  8'h00;
		ram[15'h105F] =  8'hE8;
		ram[15'h1060] =  8'h87;
		ram[15'h1061] =  8'h06;
		ram[15'h1062] =  8'h20;
		ram[15'h1063] =  8'h12;
		ram[15'h1064] =  8'hBD;
		ram[15'h1065] =  8'h9B;
		ram[15'h1066] =  8'hB6;
		ram[15'h1067] =  8'h53;
		ram[15'h1068] =  8'h72;
		ram[15'h1069] =  8'hE5;
		ram[15'h106A] =  8'hA1;
		ram[15'h106B] =  8'h51;
		ram[15'h106C] =  8'h13;
		ram[15'h106D] =  8'hBD;
		ram[15'h106E] =  8'hF1;
		ram[15'h106F] =  8'h20;
		ram[15'h1070] =  8'h00;
		ram[15'h1071] =  8'h00;
		ram[15'h1072] =  8'h00;
		ram[15'h1073] =  8'h00;
		ram[15'h1074] =  8'h00;
		ram[15'h1075] =  8'h00;
		ram[15'h1076] =  8'h00;
		ram[15'h1077] =  8'h00;
		ram[15'h1078] =  8'h00;
		ram[15'h1079] =  8'h00;
		ram[15'h107A] =  8'h00;
		ram[15'h107B] =  8'h00;
		ram[15'h107C] =  8'h00;
		ram[15'h107D] =  8'h00;
		ram[15'h107E] =  8'h00;
		ram[15'h107F] =  8'h00;
		ram[15'h1080] =  8'h00;
		ram[15'h1081] =  8'h00;
		ram[15'h1082] =  8'h00;
		ram[15'h1083] =  8'h00;
		ram[15'h1084] =  8'h00;
		ram[15'h1085] =  8'hFF;
		ram[15'h1086] =  8'hFF;
		ram[15'h1087] =  8'h00;
		ram[15'h1088] =  8'h00;
		ram[15'h1089] =  8'h00;
		ram[15'h108A] =  8'h00;
		ram[15'h108B] =  8'h00;
		ram[15'h108C] =  8'h00;
		ram[15'h108D] =  8'h00;
		ram[15'h108E] =  8'h00;
		ram[15'h108F] =  8'h00;
		ram[15'h1090] =  8'h00;
		ram[15'h1091] =  8'h00;
		ram[15'h1092] =  8'h00;
		ram[15'h1093] =  8'h00;
		ram[15'h1094] =  8'h00;
		ram[15'h1095] =  8'h00;
		ram[15'h1096] =  8'h00;
		ram[15'h1097] =  8'h22;
		ram[15'h1098] =  8'h7D;
		ram[15'h1099] =  8'hD5;
		ram[15'h109A] =  8'h25;
		ram[15'h109B] =  8'h6C;
		ram[15'h109C] =  8'h64;
		ram[15'h109D] =  8'h20;
		ram[15'h109E] =  8'h3C;
		ram[15'h109F] =  8'h69;
		ram[15'h10A0] =  8'h78;
		ram[15'h10A1] =  8'h2C;
		ram[15'h10A2] =  8'h69;
		ram[15'h10A3] =  8'h79;
		ram[15'h10A4] =  8'h3E;
		ram[15'h10A5] =  8'h2C;
		ram[15'h10A6] =  8'h6E;
		ram[15'h10A7] =  8'h6E;
		ram[15'h10A8] =  8'h6E;
		ram[15'h10A9] =  8'h6E;
		ram[15'h10AA] =  8'h2E;
		ram[15'h10AB] =  8'h2E;
		ram[15'h10AC] =  8'h2E;
		ram[15'h10AD] =  8'h2E;
		ram[15'h10AE] =  8'h2E;
		ram[15'h10AF] =  8'h2E;
		ram[15'h10B0] =  8'h2E;
		ram[15'h10B1] =  8'h2E;
		ram[15'h10B2] =  8'h2E;
		ram[15'h10B3] =  8'h2E;
		ram[15'h10B4] =  8'h2E;
		ram[15'h10B5] =  8'h2E;
		ram[15'h10B6] =  8'h2E;
		ram[15'h10B7] =  8'h2E;
		ram[15'h10B8] =  8'h2E;
		ram[15'h10B9] =  8'h24;
		ram[15'h10BA] =  8'hD7;
		ram[15'h10BB] =  8'h0A;
		ram[15'h10BC] =  8'h00;
		ram[15'h10BD] =  8'h00;
		ram[15'h10BE] =  8'h00;
		ram[15'h10BF] =  8'hA8;
		ram[15'h10C0] =  8'hB3;
		ram[15'h10C1] =  8'h2A;
		ram[15'h10C2] =  8'h1D;
		ram[15'h10C3] =  8'h8E;
		ram[15'h10C4] =  8'h7F;
		ram[15'h10C5] =  8'hAC;
		ram[15'h10C6] =  8'h42;
		ram[15'h10C7] =  8'h3A;
		ram[15'h10C8] =  8'h00;
		ram[15'h10C9] =  8'h3A;
		ram[15'h10CA] =  8'h00;
		ram[15'h10CB] =  8'hC6;
		ram[15'h10CC] =  8'hB1;
		ram[15'h10CD] =  8'h8E;
		ram[15'h10CE] =  8'hEF;
		ram[15'h10CF] =  8'h10;
		ram[15'h10D0] =  8'h00;
		ram[15'h10D1] =  8'h00;
		ram[15'h10D2] =  8'h00;
		ram[15'h10D3] =  8'h00;
		ram[15'h10D4] =  8'h00;
		ram[15'h10D5] =  8'h00;
		ram[15'h10D6] =  8'h00;
		ram[15'h10D7] =  8'h00;
		ram[15'h10D8] =  8'h00;
		ram[15'h10D9] =  8'h00;
		ram[15'h10DA] =  8'h00;
		ram[15'h10DB] =  8'h00;
		ram[15'h10DC] =  8'h00;
		ram[15'h10DD] =  8'h00;
		ram[15'h10DE] =  8'h00;
		ram[15'h10DF] =  8'h00;
		ram[15'h10E0] =  8'h00;
		ram[15'h10E1] =  8'h00;
		ram[15'h10E2] =  8'h00;
		ram[15'h10E3] =  8'h00;
		ram[15'h10E4] =  8'h00;
		ram[15'h10E5] =  8'h00;
		ram[15'h10E6] =  8'h00;
		ram[15'h10E7] =  8'hFF;
		ram[15'h10E8] =  8'h00;
		ram[15'h10E9] =  8'h00;
		ram[15'h10EA] =  8'h00;
		ram[15'h10EB] =  8'h00;
		ram[15'h10EC] =  8'h00;
		ram[15'h10ED] =  8'h00;
		ram[15'h10EE] =  8'h00;
		ram[15'h10EF] =  8'h00;
		ram[15'h10F0] =  8'h00;
		ram[15'h10F1] =  8'h00;
		ram[15'h10F2] =  8'h00;
		ram[15'h10F3] =  8'hD7;
		ram[15'h10F4] =  8'hFF;
		ram[15'h10F5] =  8'h00;
		ram[15'h10F6] =  8'h00;
		ram[15'h10F7] =  8'hB0;
		ram[15'h10F8] =  8'h81;
		ram[15'h10F9] =  8'h89;
		ram[15'h10FA] =  8'h35;
		ram[15'h10FB] =  8'h6C;
		ram[15'h10FC] =  8'h64;
		ram[15'h10FD] =  8'h20;
		ram[15'h10FE] =  8'h61;
		ram[15'h10FF] =  8'h2C;
		ram[15'h1100] =  8'h3C;
		ram[15'h1101] =  8'h28;
		ram[15'h1102] =  8'h62;
		ram[15'h1103] =  8'h63;
		ram[15'h1104] =  8'h29;
		ram[15'h1105] =  8'h2C;
		ram[15'h1106] =  8'h28;
		ram[15'h1107] =  8'h64;
		ram[15'h1108] =  8'h65;
		ram[15'h1109] =  8'h29;
		ram[15'h110A] =  8'h3E;
		ram[15'h110B] =  8'h2E;
		ram[15'h110C] =  8'h2E;
		ram[15'h110D] =  8'h2E;
		ram[15'h110E] =  8'h2E;
		ram[15'h110F] =  8'h2E;
		ram[15'h1110] =  8'h2E;
		ram[15'h1111] =  8'h2E;
		ram[15'h1112] =  8'h2E;
		ram[15'h1113] =  8'h2E;
		ram[15'h1114] =  8'h2E;
		ram[15'h1115] =  8'h2E;
		ram[15'h1116] =  8'h2E;
		ram[15'h1117] =  8'h2E;
		ram[15'h1118] =  8'h2E;
		ram[15'h1119] =  8'h24;
		ram[15'h111A] =  8'hD7;
		ram[15'h111B] =  8'h06;
		ram[15'h111C] =  8'h00;
		ram[15'h111D] =  8'h00;
		ram[15'h111E] =  8'h00;
		ram[15'h111F] =  8'h07;
		ram[15'h1120] =  8'hC4;
		ram[15'h1121] =  8'h9D;
		ram[15'h1122] =  8'hF4;
		ram[15'h1123] =  8'h3D;
		ram[15'h1124] =  8'hD1;
		ram[15'h1125] =  8'h39;
		ram[15'h1126] =  8'h03;
		ram[15'h1127] =  8'h89;
		ram[15'h1128] =  8'hDE;
		ram[15'h1129] =  8'h55;
		ram[15'h112A] =  8'h74;
		ram[15'h112B] =  8'h53;
		ram[15'h112C] =  8'hC0;
		ram[15'h112D] =  8'h09;
		ram[15'h112E] =  8'h55;
		ram[15'h112F] =  8'h38;
		ram[15'h1130] =  8'h00;
		ram[15'h1131] =  8'h00;
		ram[15'h1132] =  8'h00;
		ram[15'h1133] =  8'h00;
		ram[15'h1134] =  8'h00;
		ram[15'h1135] =  8'h00;
		ram[15'h1136] =  8'h00;
		ram[15'h1137] =  8'h00;
		ram[15'h1138] =  8'h00;
		ram[15'h1139] =  8'h00;
		ram[15'h113A] =  8'h00;
		ram[15'h113B] =  8'h00;
		ram[15'h113C] =  8'h00;
		ram[15'h113D] =  8'h00;
		ram[15'h113E] =  8'h00;
		ram[15'h113F] =  8'h00;
		ram[15'h1140] =  8'h00;
		ram[15'h1141] =  8'h00;
		ram[15'h1142] =  8'h00;
		ram[15'h1143] =  8'h00;
		ram[15'h1144] =  8'h00;
		ram[15'h1145] =  8'h00;
		ram[15'h1146] =  8'h00;
		ram[15'h1147] =  8'h00;
		ram[15'h1148] =  8'h00;
		ram[15'h1149] =  8'h00;
		ram[15'h114A] =  8'h00;
		ram[15'h114B] =  8'h00;
		ram[15'h114C] =  8'h00;
		ram[15'h114D] =  8'h00;
		ram[15'h114E] =  8'h00;
		ram[15'h114F] =  8'h00;
		ram[15'h1150] =  8'h00;
		ram[15'h1151] =  8'h00;
		ram[15'h1152] =  8'h00;
		ram[15'h1153] =  8'h00;
		ram[15'h1154] =  8'hFF;
		ram[15'h1155] =  8'h00;
		ram[15'h1156] =  8'h00;
		ram[15'h1157] =  8'hF1;
		ram[15'h1158] =  8'hDA;
		ram[15'h1159] =  8'hB5;
		ram[15'h115A] =  8'h56;
		ram[15'h115B] =  8'h6C;
		ram[15'h115C] =  8'h64;
		ram[15'h115D] =  8'h20;
		ram[15'h115E] =  8'h3C;
		ram[15'h115F] =  8'h62;
		ram[15'h1160] =  8'h2C;
		ram[15'h1161] =  8'h63;
		ram[15'h1162] =  8'h2C;
		ram[15'h1163] =  8'h64;
		ram[15'h1164] =  8'h2C;
		ram[15'h1165] =  8'h65;
		ram[15'h1166] =  8'h2C;
		ram[15'h1167] =  8'h68;
		ram[15'h1168] =  8'h2C;
		ram[15'h1169] =  8'h6C;
		ram[15'h116A] =  8'h2C;
		ram[15'h116B] =  8'h28;
		ram[15'h116C] =  8'h68;
		ram[15'h116D] =  8'h6C;
		ram[15'h116E] =  8'h29;
		ram[15'h116F] =  8'h2C;
		ram[15'h1170] =  8'h61;
		ram[15'h1171] =  8'h3E;
		ram[15'h1172] =  8'h2C;
		ram[15'h1173] =  8'h6E;
		ram[15'h1174] =  8'h6E;
		ram[15'h1175] =  8'h2E;
		ram[15'h1176] =  8'h2E;
		ram[15'h1177] =  8'h2E;
		ram[15'h1178] =  8'h2E;
		ram[15'h1179] =  8'h24;
		ram[15'h117A] =  8'hD7;
		ram[15'h117B] =  8'hDD;
		ram[15'h117C] =  8'h36;
		ram[15'h117D] =  8'h01;
		ram[15'h117E] =  8'h00;
		ram[15'h117F] =  8'h45;
		ram[15'h1180] =  8'h1B;
		ram[15'h1181] =  8'h39;
		ram[15'h1182] =  8'h00;
		ram[15'h1183] =  8'h39;
		ram[15'h1184] =  8'h00;
		ram[15'h1185] =  8'hC1;
		ram[15'h1186] =  8'hD5;
		ram[15'h1187] =  8'hC7;
		ram[15'h1188] =  8'h61;
		ram[15'h1189] =  8'hC4;
		ram[15'h118A] =  8'hBD;
		ram[15'h118B] =  8'hC0;
		ram[15'h118C] =  8'h85;
		ram[15'h118D] =  8'h16;
		ram[15'h118E] =  8'hCD;
		ram[15'h118F] =  8'h20;
		ram[15'h1190] =  8'h00;
		ram[15'h1191] =  8'h00;
		ram[15'h1192] =  8'h00;
		ram[15'h1193] =  8'h00;
		ram[15'h1194] =  8'h00;
		ram[15'h1195] =  8'h00;
		ram[15'h1196] =  8'h00;
		ram[15'h1197] =  8'h00;
		ram[15'h1198] =  8'h00;
		ram[15'h1199] =  8'h00;
		ram[15'h119A] =  8'h00;
		ram[15'h119B] =  8'h00;
		ram[15'h119C] =  8'h00;
		ram[15'h119D] =  8'h00;
		ram[15'h119E] =  8'h00;
		ram[15'h119F] =  8'h00;
		ram[15'h11A0] =  8'h00;
		ram[15'h11A1] =  8'h00;
		ram[15'h11A2] =  8'h00;
		ram[15'h11A3] =  8'h00;
		ram[15'h11A4] =  8'h00;
		ram[15'h11A5] =  8'h00;
		ram[15'h11A6] =  8'hFF;
		ram[15'h11A7] =  8'h00;
		ram[15'h11A8] =  8'h00;
		ram[15'h11A9] =  8'h00;
		ram[15'h11AA] =  8'h00;
		ram[15'h11AB] =  8'h00;
		ram[15'h11AC] =  8'h00;
		ram[15'h11AD] =  8'h00;
		ram[15'h11AE] =  8'h00;
		ram[15'h11AF] =  8'h00;
		ram[15'h11B0] =  8'h00;
		ram[15'h11B1] =  8'h00;
		ram[15'h11B2] =  8'h00;
		ram[15'h11B3] =  8'h00;
		ram[15'h11B4] =  8'hFF;
		ram[15'h11B5] =  8'h00;
		ram[15'h11B6] =  8'h00;
		ram[15'h11B7] =  8'h26;
		ram[15'h11B8] =  8'hDB;
		ram[15'h11B9] =  8'h47;
		ram[15'h11BA] =  8'h7E;
		ram[15'h11BB] =  8'h6C;
		ram[15'h11BC] =  8'h64;
		ram[15'h11BD] =  8'h20;
		ram[15'h11BE] =  8'h28;
		ram[15'h11BF] =  8'h3C;
		ram[15'h11C0] =  8'h69;
		ram[15'h11C1] =  8'h78;
		ram[15'h11C2] =  8'h2C;
		ram[15'h11C3] =  8'h69;
		ram[15'h11C4] =  8'h79;
		ram[15'h11C5] =  8'h3E;
		ram[15'h11C6] =  8'h2B;
		ram[15'h11C7] =  8'h31;
		ram[15'h11C8] =  8'h29;
		ram[15'h11C9] =  8'h2C;
		ram[15'h11CA] =  8'h6E;
		ram[15'h11CB] =  8'h6E;
		ram[15'h11CC] =  8'h2E;
		ram[15'h11CD] =  8'h2E;
		ram[15'h11CE] =  8'h2E;
		ram[15'h11CF] =  8'h2E;
		ram[15'h11D0] =  8'h2E;
		ram[15'h11D1] =  8'h2E;
		ram[15'h11D2] =  8'h2E;
		ram[15'h11D3] =  8'h2E;
		ram[15'h11D4] =  8'h2E;
		ram[15'h11D5] =  8'h2E;
		ram[15'h11D6] =  8'h2E;
		ram[15'h11D7] =  8'h2E;
		ram[15'h11D8] =  8'h2E;
		ram[15'h11D9] =  8'h24;
		ram[15'h11DA] =  8'hD7;
		ram[15'h11DB] =  8'hDD;
		ram[15'h11DC] =  8'h46;
		ram[15'h11DD] =  8'h01;
		ram[15'h11DE] =  8'h00;
		ram[15'h11DF] =  8'h16;
		ram[15'h11E0] =  8'hD0;
		ram[15'h11E1] =  8'h39;
		ram[15'h11E2] =  8'h00;
		ram[15'h11E3] =  8'h39;
		ram[15'h11E4] =  8'h00;
		ram[15'h11E5] =  8'h60;
		ram[15'h11E6] =  8'h42;
		ram[15'h11E7] =  8'h39;
		ram[15'h11E8] =  8'h7F;
		ram[15'h11E9] =  8'h04;
		ram[15'h11EA] =  8'h04;
		ram[15'h11EB] =  8'h97;
		ram[15'h11EC] =  8'h4A;
		ram[15'h11ED] =  8'h85;
		ram[15'h11EE] =  8'hD0;
		ram[15'h11EF] =  8'h20;
		ram[15'h11F0] =  8'h18;
		ram[15'h11F1] =  8'h00;
		ram[15'h11F2] =  8'h00;
		ram[15'h11F3] =  8'h00;
		ram[15'h11F4] =  8'h00;
		ram[15'h11F5] =  8'h01;
		ram[15'h11F6] =  8'h00;
		ram[15'h11F7] =  8'h01;
		ram[15'h11F8] =  8'h00;
		ram[15'h11F9] =  8'h00;
		ram[15'h11FA] =  8'h00;
		ram[15'h11FB] =  8'h00;
		ram[15'h11FC] =  8'h00;
		ram[15'h11FD] =  8'h00;
		ram[15'h11FE] =  8'h00;
		ram[15'h11FF] =  8'h00;
		ram[15'h1200] =  8'h00;
		ram[15'h1201] =  8'h00;
		ram[15'h1202] =  8'h00;
		ram[15'h1203] =  8'h00;
		ram[15'h1204] =  8'h00;
		ram[15'h1205] =  8'h00;
		ram[15'h1206] =  8'h00;
		ram[15'h1207] =  8'hFF;
		ram[15'h1208] =  8'hFF;
		ram[15'h1209] =  8'h00;
		ram[15'h120A] =  8'h00;
		ram[15'h120B] =  8'h00;
		ram[15'h120C] =  8'h00;
		ram[15'h120D] =  8'h00;
		ram[15'h120E] =  8'h00;
		ram[15'h120F] =  8'h00;
		ram[15'h1210] =  8'h00;
		ram[15'h1211] =  8'h00;
		ram[15'h1212] =  8'h00;
		ram[15'h1213] =  8'h00;
		ram[15'h1214] =  8'h00;
		ram[15'h1215] =  8'h00;
		ram[15'h1216] =  8'h00;
		ram[15'h1217] =  8'hCC;
		ram[15'h1218] =  8'h11;
		ram[15'h1219] =  8'h06;
		ram[15'h121A] =  8'hA8;
		ram[15'h121B] =  8'h6C;
		ram[15'h121C] =  8'h64;
		ram[15'h121D] =  8'h20;
		ram[15'h121E] =  8'h3C;
		ram[15'h121F] =  8'h62;
		ram[15'h1220] =  8'h2C;
		ram[15'h1221] =  8'h63;
		ram[15'h1222] =  8'h2C;
		ram[15'h1223] =  8'h64;
		ram[15'h1224] =  8'h2C;
		ram[15'h1225] =  8'h65;
		ram[15'h1226] =  8'h3E;
		ram[15'h1227] =  8'h2C;
		ram[15'h1228] =  8'h28;
		ram[15'h1229] =  8'h3C;
		ram[15'h122A] =  8'h69;
		ram[15'h122B] =  8'h78;
		ram[15'h122C] =  8'h2C;
		ram[15'h122D] =  8'h69;
		ram[15'h122E] =  8'h79;
		ram[15'h122F] =  8'h3E;
		ram[15'h1230] =  8'h2B;
		ram[15'h1231] =  8'h31;
		ram[15'h1232] =  8'h29;
		ram[15'h1233] =  8'h2E;
		ram[15'h1234] =  8'h2E;
		ram[15'h1235] =  8'h2E;
		ram[15'h1236] =  8'h2E;
		ram[15'h1237] =  8'h2E;
		ram[15'h1238] =  8'h2E;
		ram[15'h1239] =  8'h24;
		ram[15'h123A] =  8'hD7;
		ram[15'h123B] =  8'hDD;
		ram[15'h123C] =  8'h66;
		ram[15'h123D] =  8'h01;
		ram[15'h123E] =  8'h00;
		ram[15'h123F] =  8'hE0;
		ram[15'h1240] =  8'h84;
		ram[15'h1241] =  8'h39;
		ram[15'h1242] =  8'h00;
		ram[15'h1243] =  8'h39;
		ram[15'h1244] =  8'h00;
		ram[15'h1245] =  8'h52;
		ram[15'h1246] =  8'h9C;
		ram[15'h1247] =  8'h99;
		ram[15'h1248] =  8'hA7;
		ram[15'h1249] =  8'hB6;
		ram[15'h124A] =  8'h49;
		ram[15'h124B] =  8'h93;
		ram[15'h124C] =  8'h00;
		ram[15'h124D] =  8'hAD;
		ram[15'h124E] =  8'hEE;
		ram[15'h124F] =  8'h20;
		ram[15'h1250] =  8'h08;
		ram[15'h1251] =  8'h00;
		ram[15'h1252] =  8'h00;
		ram[15'h1253] =  8'h00;
		ram[15'h1254] =  8'h00;
		ram[15'h1255] =  8'h01;
		ram[15'h1256] =  8'h00;
		ram[15'h1257] =  8'h01;
		ram[15'h1258] =  8'h00;
		ram[15'h1259] =  8'h00;
		ram[15'h125A] =  8'h00;
		ram[15'h125B] =  8'h00;
		ram[15'h125C] =  8'h00;
		ram[15'h125D] =  8'h00;
		ram[15'h125E] =  8'h00;
		ram[15'h125F] =  8'h00;
		ram[15'h1260] =  8'h00;
		ram[15'h1261] =  8'h00;
		ram[15'h1262] =  8'h00;
		ram[15'h1263] =  8'h00;
		ram[15'h1264] =  8'h00;
		ram[15'h1265] =  8'h00;
		ram[15'h1266] =  8'h00;
		ram[15'h1267] =  8'hFF;
		ram[15'h1268] =  8'hFF;
		ram[15'h1269] =  8'h00;
		ram[15'h126A] =  8'h00;
		ram[15'h126B] =  8'h00;
		ram[15'h126C] =  8'h00;
		ram[15'h126D] =  8'h00;
		ram[15'h126E] =  8'h00;
		ram[15'h126F] =  8'h00;
		ram[15'h1270] =  8'h00;
		ram[15'h1271] =  8'h00;
		ram[15'h1272] =  8'h00;
		ram[15'h1273] =  8'h00;
		ram[15'h1274] =  8'h00;
		ram[15'h1275] =  8'h00;
		ram[15'h1276] =  8'h00;
		ram[15'h1277] =  8'hFA;
		ram[15'h1278] =  8'h2A;
		ram[15'h1279] =  8'h4D;
		ram[15'h127A] =  8'h03;
		ram[15'h127B] =  8'h6C;
		ram[15'h127C] =  8'h64;
		ram[15'h127D] =  8'h20;
		ram[15'h127E] =  8'h3C;
		ram[15'h127F] =  8'h68;
		ram[15'h1280] =  8'h2C;
		ram[15'h1281] =  8'h6C;
		ram[15'h1282] =  8'h3E;
		ram[15'h1283] =  8'h2C;
		ram[15'h1284] =  8'h28;
		ram[15'h1285] =  8'h3C;
		ram[15'h1286] =  8'h69;
		ram[15'h1287] =  8'h78;
		ram[15'h1288] =  8'h2C;
		ram[15'h1289] =  8'h69;
		ram[15'h128A] =  8'h79;
		ram[15'h128B] =  8'h3E;
		ram[15'h128C] =  8'h2B;
		ram[15'h128D] =  8'h31;
		ram[15'h128E] =  8'h29;
		ram[15'h128F] =  8'h2E;
		ram[15'h1290] =  8'h2E;
		ram[15'h1291] =  8'h2E;
		ram[15'h1292] =  8'h2E;
		ram[15'h1293] =  8'h2E;
		ram[15'h1294] =  8'h2E;
		ram[15'h1295] =  8'h2E;
		ram[15'h1296] =  8'h2E;
		ram[15'h1297] =  8'h2E;
		ram[15'h1298] =  8'h2E;
		ram[15'h1299] =  8'h24;
		ram[15'h129A] =  8'hD7;
		ram[15'h129B] =  8'hDD;
		ram[15'h129C] =  8'h7E;
		ram[15'h129D] =  8'h01;
		ram[15'h129E] =  8'h00;
		ram[15'h129F] =  8'hB6;
		ram[15'h12A0] =  8'hD8;
		ram[15'h12A1] =  8'h39;
		ram[15'h12A2] =  8'h00;
		ram[15'h12A3] =  8'h39;
		ram[15'h12A4] =  8'h00;
		ram[15'h12A5] =  8'h12;
		ram[15'h12A6] =  8'hC6;
		ram[15'h12A7] =  8'h07;
		ram[15'h12A8] =  8'hDF;
		ram[15'h12A9] =  8'hD0;
		ram[15'h12AA] =  8'h9C;
		ram[15'h12AB] =  8'h43;
		ram[15'h12AC] =  8'hA6;
		ram[15'h12AD] =  8'hE5;
		ram[15'h12AE] =  8'hA0;
		ram[15'h12AF] =  8'h20;
		ram[15'h12B0] =  8'h00;
		ram[15'h12B1] =  8'h00;
		ram[15'h12B2] =  8'h00;
		ram[15'h12B3] =  8'h00;
		ram[15'h12B4] =  8'h00;
		ram[15'h12B5] =  8'h01;
		ram[15'h12B6] =  8'h00;
		ram[15'h12B7] =  8'h01;
		ram[15'h12B8] =  8'h00;
		ram[15'h12B9] =  8'h00;
		ram[15'h12BA] =  8'h00;
		ram[15'h12BB] =  8'h00;
		ram[15'h12BC] =  8'h00;
		ram[15'h12BD] =  8'h00;
		ram[15'h12BE] =  8'h00;
		ram[15'h12BF] =  8'h00;
		ram[15'h12C0] =  8'h00;
		ram[15'h12C1] =  8'h00;
		ram[15'h12C2] =  8'h00;
		ram[15'h12C3] =  8'h00;
		ram[15'h12C4] =  8'h00;
		ram[15'h12C5] =  8'h00;
		ram[15'h12C6] =  8'h00;
		ram[15'h12C7] =  8'hFF;
		ram[15'h12C8] =  8'hFF;
		ram[15'h12C9] =  8'h00;
		ram[15'h12CA] =  8'h00;
		ram[15'h12CB] =  8'h00;
		ram[15'h12CC] =  8'h00;
		ram[15'h12CD] =  8'h00;
		ram[15'h12CE] =  8'h00;
		ram[15'h12CF] =  8'h00;
		ram[15'h12D0] =  8'h00;
		ram[15'h12D1] =  8'h00;
		ram[15'h12D2] =  8'h00;
		ram[15'h12D3] =  8'h00;
		ram[15'h12D4] =  8'h00;
		ram[15'h12D5] =  8'h00;
		ram[15'h12D6] =  8'h00;
		ram[15'h12D7] =  8'hA5;
		ram[15'h12D8] =  8'hE9;
		ram[15'h12D9] =  8'hAC;
		ram[15'h12DA] =  8'h64;
		ram[15'h12DB] =  8'h6C;
		ram[15'h12DC] =  8'h64;
		ram[15'h12DD] =  8'h20;
		ram[15'h12DE] =  8'h61;
		ram[15'h12DF] =  8'h2C;
		ram[15'h12E0] =  8'h28;
		ram[15'h12E1] =  8'h3C;
		ram[15'h12E2] =  8'h69;
		ram[15'h12E3] =  8'h78;
		ram[15'h12E4] =  8'h2C;
		ram[15'h12E5] =  8'h69;
		ram[15'h12E6] =  8'h79;
		ram[15'h12E7] =  8'h3E;
		ram[15'h12E8] =  8'h2B;
		ram[15'h12E9] =  8'h31;
		ram[15'h12EA] =  8'h29;
		ram[15'h12EB] =  8'h2E;
		ram[15'h12EC] =  8'h2E;
		ram[15'h12ED] =  8'h2E;
		ram[15'h12EE] =  8'h2E;
		ram[15'h12EF] =  8'h2E;
		ram[15'h12F0] =  8'h2E;
		ram[15'h12F1] =  8'h2E;
		ram[15'h12F2] =  8'h2E;
		ram[15'h12F3] =  8'h2E;
		ram[15'h12F4] =  8'h2E;
		ram[15'h12F5] =  8'h2E;
		ram[15'h12F6] =  8'h2E;
		ram[15'h12F7] =  8'h2E;
		ram[15'h12F8] =  8'h2E;
		ram[15'h12F9] =  8'h24;
		ram[15'h12FA] =  8'hD7;
		ram[15'h12FB] =  8'hDD;
		ram[15'h12FC] =  8'h26;
		ram[15'h12FD] =  8'h00;
		ram[15'h12FE] =  8'h00;
		ram[15'h12FF] =  8'h53;
		ram[15'h1300] =  8'h3C;
		ram[15'h1301] =  8'h40;
		ram[15'h1302] =  8'h46;
		ram[15'h1303] =  8'h79;
		ram[15'h1304] =  8'hE1;
		ram[15'h1305] =  8'h11;
		ram[15'h1306] =  8'h77;
		ram[15'h1307] =  8'h07;
		ram[15'h1308] =  8'hC1;
		ram[15'h1309] =  8'hFA;
		ram[15'h130A] =  8'h1A;
		ram[15'h130B] =  8'h81;
		ram[15'h130C] =  8'hAD;
		ram[15'h130D] =  8'h9B;
		ram[15'h130E] =  8'h5D;
		ram[15'h130F] =  8'h20;
		ram[15'h1310] =  8'h08;
		ram[15'h1311] =  8'h00;
		ram[15'h1312] =  8'h00;
		ram[15'h1313] =  8'h00;
		ram[15'h1314] =  8'h00;
		ram[15'h1315] =  8'h00;
		ram[15'h1316] =  8'h00;
		ram[15'h1317] =  8'h00;
		ram[15'h1318] =  8'h00;
		ram[15'h1319] =  8'h00;
		ram[15'h131A] =  8'h00;
		ram[15'h131B] =  8'h00;
		ram[15'h131C] =  8'h00;
		ram[15'h131D] =  8'h00;
		ram[15'h131E] =  8'h00;
		ram[15'h131F] =  8'h00;
		ram[15'h1320] =  8'h00;
		ram[15'h1321] =  8'h00;
		ram[15'h1322] =  8'h00;
		ram[15'h1323] =  8'h00;
		ram[15'h1324] =  8'h00;
		ram[15'h1325] =  8'h00;
		ram[15'h1326] =  8'h00;
		ram[15'h1327] =  8'h00;
		ram[15'h1328] =  8'h00;
		ram[15'h1329] =  8'h00;
		ram[15'h132A] =  8'h00;
		ram[15'h132B] =  8'h00;
		ram[15'h132C] =  8'h00;
		ram[15'h132D] =  8'h00;
		ram[15'h132E] =  8'h00;
		ram[15'h132F] =  8'h00;
		ram[15'h1330] =  8'h00;
		ram[15'h1331] =  8'h00;
		ram[15'h1332] =  8'h00;
		ram[15'h1333] =  8'h00;
		ram[15'h1334] =  8'hFF;
		ram[15'h1335] =  8'h00;
		ram[15'h1336] =  8'h00;
		ram[15'h1337] =  8'h24;
		ram[15'h1338] =  8'hE8;
		ram[15'h1339] =  8'h82;
		ram[15'h133A] =  8'h8B;
		ram[15'h133B] =  8'h6C;
		ram[15'h133C] =  8'h64;
		ram[15'h133D] =  8'h20;
		ram[15'h133E] =  8'h3C;
		ram[15'h133F] =  8'h69;
		ram[15'h1340] =  8'h78;
		ram[15'h1341] =  8'h68;
		ram[15'h1342] =  8'h2C;
		ram[15'h1343] =  8'h69;
		ram[15'h1344] =  8'h78;
		ram[15'h1345] =  8'h6C;
		ram[15'h1346] =  8'h2C;
		ram[15'h1347] =  8'h69;
		ram[15'h1348] =  8'h79;
		ram[15'h1349] =  8'h68;
		ram[15'h134A] =  8'h2C;
		ram[15'h134B] =  8'h69;
		ram[15'h134C] =  8'h79;
		ram[15'h134D] =  8'h6C;
		ram[15'h134E] =  8'h3E;
		ram[15'h134F] =  8'h2C;
		ram[15'h1350] =  8'h6E;
		ram[15'h1351] =  8'h6E;
		ram[15'h1352] =  8'h2E;
		ram[15'h1353] =  8'h2E;
		ram[15'h1354] =  8'h2E;
		ram[15'h1355] =  8'h2E;
		ram[15'h1356] =  8'h2E;
		ram[15'h1357] =  8'h2E;
		ram[15'h1358] =  8'h2E;
		ram[15'h1359] =  8'h24;
		ram[15'h135A] =  8'hD7;
		ram[15'h135B] =  8'h40;
		ram[15'h135C] =  8'h00;
		ram[15'h135D] =  8'h00;
		ram[15'h135E] =  8'h00;
		ram[15'h135F] =  8'hA4;
		ram[15'h1360] =  8'h72;
		ram[15'h1361] =  8'h24;
		ram[15'h1362] =  8'hA0;
		ram[15'h1363] =  8'hAC;
		ram[15'h1364] =  8'h61;
		ram[15'h1365] =  8'h3A;
		ram[15'h1366] =  8'h00;
		ram[15'h1367] =  8'hC7;
		ram[15'h1368] =  8'h82;
		ram[15'h1369] =  8'h8F;
		ram[15'h136A] =  8'h71;
		ram[15'h136B] =  8'h97;
		ram[15'h136C] =  8'h8F;
		ram[15'h136D] =  8'h8E;
		ram[15'h136E] =  8'hEF;
		ram[15'h136F] =  8'h3F;
		ram[15'h1370] =  8'h00;
		ram[15'h1371] =  8'h00;
		ram[15'h1372] =  8'h00;
		ram[15'h1373] =  8'h00;
		ram[15'h1374] =  8'h00;
		ram[15'h1375] =  8'h00;
		ram[15'h1376] =  8'h00;
		ram[15'h1377] =  8'h00;
		ram[15'h1378] =  8'h00;
		ram[15'h1379] =  8'h00;
		ram[15'h137A] =  8'h00;
		ram[15'h137B] =  8'h00;
		ram[15'h137C] =  8'h00;
		ram[15'h137D] =  8'h00;
		ram[15'h137E] =  8'h00;
		ram[15'h137F] =  8'h00;
		ram[15'h1380] =  8'h00;
		ram[15'h1381] =  8'h00;
		ram[15'h1382] =  8'h00;
		ram[15'h1383] =  8'h00;
		ram[15'h1384] =  8'h00;
		ram[15'h1385] =  8'h00;
		ram[15'h1386] =  8'h00;
		ram[15'h1387] =  8'hFF;
		ram[15'h1388] =  8'h00;
		ram[15'h1389] =  8'h00;
		ram[15'h138A] =  8'h00;
		ram[15'h138B] =  8'h00;
		ram[15'h138C] =  8'h00;
		ram[15'h138D] =  8'h00;
		ram[15'h138E] =  8'h00;
		ram[15'h138F] =  8'hFF;
		ram[15'h1390] =  8'hFF;
		ram[15'h1391] =  8'hFF;
		ram[15'h1392] =  8'hFF;
		ram[15'h1393] =  8'hD7;
		ram[15'h1394] =  8'hFF;
		ram[15'h1395] =  8'h00;
		ram[15'h1396] =  8'h00;
		ram[15'h1397] =  8'h74;
		ram[15'h1398] =  8'h4B;
		ram[15'h1399] =  8'h01;
		ram[15'h139A] =  8'h18;
		ram[15'h139B] =  8'h6C;
		ram[15'h139C] =  8'h64;
		ram[15'h139D] =  8'h20;
		ram[15'h139E] =  8'h3C;
		ram[15'h139F] =  8'h62;
		ram[15'h13A0] =  8'h63;
		ram[15'h13A1] =  8'h64;
		ram[15'h13A2] =  8'h65;
		ram[15'h13A3] =  8'h68;
		ram[15'h13A4] =  8'h6C;
		ram[15'h13A5] =  8'h61;
		ram[15'h13A6] =  8'h3E;
		ram[15'h13A7] =  8'h2C;
		ram[15'h13A8] =  8'h3C;
		ram[15'h13A9] =  8'h62;
		ram[15'h13AA] =  8'h63;
		ram[15'h13AB] =  8'h64;
		ram[15'h13AC] =  8'h65;
		ram[15'h13AD] =  8'h68;
		ram[15'h13AE] =  8'h6C;
		ram[15'h13AF] =  8'h61;
		ram[15'h13B0] =  8'h3E;
		ram[15'h13B1] =  8'h2E;
		ram[15'h13B2] =  8'h2E;
		ram[15'h13B3] =  8'h2E;
		ram[15'h13B4] =  8'h2E;
		ram[15'h13B5] =  8'h2E;
		ram[15'h13B6] =  8'h2E;
		ram[15'h13B7] =  8'h2E;
		ram[15'h13B8] =  8'h2E;
		ram[15'h13B9] =  8'h24;
		ram[15'h13BA] =  8'hD7;
		ram[15'h13BB] =  8'hDD;
		ram[15'h13BC] =  8'h40;
		ram[15'h13BD] =  8'h00;
		ram[15'h13BE] =  8'h00;
		ram[15'h13BF] =  8'hC5;
		ram[15'h13C0] =  8'hBC;
		ram[15'h13C1] =  8'h3A;
		ram[15'h13C2] =  8'h00;
		ram[15'h13C3] =  8'h3A;
		ram[15'h13C4] =  8'h00;
		ram[15'h13C5] =  8'h3A;
		ram[15'h13C6] =  8'h00;
		ram[15'h13C7] =  8'hC2;
		ram[15'h13C8] =  8'h2F;
		ram[15'h13C9] =  8'hC0;
		ram[15'h13CA] =  8'h98;
		ram[15'h13CB] =  8'h83;
		ram[15'h13CC] =  8'h1F;
		ram[15'h13CD] =  8'hCD;
		ram[15'h13CE] =  8'h3B;
		ram[15'h13CF] =  8'h20;
		ram[15'h13D0] =  8'h3F;
		ram[15'h13D1] =  8'h00;
		ram[15'h13D2] =  8'h00;
		ram[15'h13D3] =  8'h00;
		ram[15'h13D4] =  8'h00;
		ram[15'h13D5] =  8'h00;
		ram[15'h13D6] =  8'h00;
		ram[15'h13D7] =  8'h00;
		ram[15'h13D8] =  8'h00;
		ram[15'h13D9] =  8'h00;
		ram[15'h13DA] =  8'h00;
		ram[15'h13DB] =  8'h00;
		ram[15'h13DC] =  8'h00;
		ram[15'h13DD] =  8'h00;
		ram[15'h13DE] =  8'h00;
		ram[15'h13DF] =  8'h00;
		ram[15'h13E0] =  8'h00;
		ram[15'h13E1] =  8'h00;
		ram[15'h13E2] =  8'h00;
		ram[15'h13E3] =  8'h00;
		ram[15'h13E4] =  8'h00;
		ram[15'h13E5] =  8'h00;
		ram[15'h13E6] =  8'h00;
		ram[15'h13E7] =  8'hFF;
		ram[15'h13E8] =  8'h00;
		ram[15'h13E9] =  8'h00;
		ram[15'h13EA] =  8'h00;
		ram[15'h13EB] =  8'h00;
		ram[15'h13EC] =  8'h00;
		ram[15'h13ED] =  8'h00;
		ram[15'h13EE] =  8'h00;
		ram[15'h13EF] =  8'hFF;
		ram[15'h13F0] =  8'hFF;
		ram[15'h13F1] =  8'hFF;
		ram[15'h13F2] =  8'hFF;
		ram[15'h13F3] =  8'hD7;
		ram[15'h13F4] =  8'hFF;
		ram[15'h13F5] =  8'h00;
		ram[15'h13F6] =  8'h00;
		ram[15'h13F7] =  8'h47;
		ram[15'h13F8] =  8'h8B;
		ram[15'h13F9] =  8'hA3;
		ram[15'h13FA] =  8'h6B;
		ram[15'h13FB] =  8'h6C;
		ram[15'h13FC] =  8'h64;
		ram[15'h13FD] =  8'h20;
		ram[15'h13FE] =  8'h3C;
		ram[15'h13FF] =  8'h62;
		ram[15'h1400] =  8'h63;
		ram[15'h1401] =  8'h64;
		ram[15'h1402] =  8'h65;
		ram[15'h1403] =  8'h78;
		ram[15'h1404] =  8'h79;
		ram[15'h1405] =  8'h61;
		ram[15'h1406] =  8'h3E;
		ram[15'h1407] =  8'h2C;
		ram[15'h1408] =  8'h3C;
		ram[15'h1409] =  8'h62;
		ram[15'h140A] =  8'h63;
		ram[15'h140B] =  8'h64;
		ram[15'h140C] =  8'h65;
		ram[15'h140D] =  8'h78;
		ram[15'h140E] =  8'h79;
		ram[15'h140F] =  8'h61;
		ram[15'h1410] =  8'h3E;
		ram[15'h1411] =  8'h2E;
		ram[15'h1412] =  8'h2E;
		ram[15'h1413] =  8'h2E;
		ram[15'h1414] =  8'h2E;
		ram[15'h1415] =  8'h2E;
		ram[15'h1416] =  8'h2E;
		ram[15'h1417] =  8'h2E;
		ram[15'h1418] =  8'h2E;
		ram[15'h1419] =  8'h24;
		ram[15'h141A] =  8'hD7;
		ram[15'h141B] =  8'h32;
		ram[15'h141C] =  8'h3A;
		ram[15'h141D] =  8'h00;
		ram[15'h141E] =  8'h00;
		ram[15'h141F] =  8'h68;
		ram[15'h1420] =  8'hFD;
		ram[15'h1421] =  8'hEC;
		ram[15'h1422] =  8'hF4;
		ram[15'h1423] =  8'hA0;
		ram[15'h1424] =  8'h44;
		ram[15'h1425] =  8'h43;
		ram[15'h1426] =  8'hB5;
		ram[15'h1427] =  8'h53;
		ram[15'h1428] =  8'h06;
		ram[15'h1429] =  8'hBA;
		ram[15'h142A] =  8'hCD;
		ram[15'h142B] =  8'hD2;
		ram[15'h142C] =  8'h4F;
		ram[15'h142D] =  8'hD8;
		ram[15'h142E] =  8'h1F;
		ram[15'h142F] =  8'h08;
		ram[15'h1430] =  8'h00;
		ram[15'h1431] =  8'h00;
		ram[15'h1432] =  8'h00;
		ram[15'h1433] =  8'h00;
		ram[15'h1434] =  8'h00;
		ram[15'h1435] =  8'h00;
		ram[15'h1436] =  8'h00;
		ram[15'h1437] =  8'h00;
		ram[15'h1438] =  8'h00;
		ram[15'h1439] =  8'h00;
		ram[15'h143A] =  8'h00;
		ram[15'h143B] =  8'h00;
		ram[15'h143C] =  8'h00;
		ram[15'h143D] =  8'h00;
		ram[15'h143E] =  8'h00;
		ram[15'h143F] =  8'h00;
		ram[15'h1440] =  8'h00;
		ram[15'h1441] =  8'h00;
		ram[15'h1442] =  8'h00;
		ram[15'h1443] =  8'h00;
		ram[15'h1444] =  8'h00;
		ram[15'h1445] =  8'h00;
		ram[15'h1446] =  8'h00;
		ram[15'h1447] =  8'hFF;
		ram[15'h1448] =  8'h00;
		ram[15'h1449] =  8'h00;
		ram[15'h144A] =  8'h00;
		ram[15'h144B] =  8'h00;
		ram[15'h144C] =  8'h00;
		ram[15'h144D] =  8'h00;
		ram[15'h144E] =  8'h00;
		ram[15'h144F] =  8'h00;
		ram[15'h1450] =  8'h00;
		ram[15'h1451] =  8'h00;
		ram[15'h1452] =  8'h00;
		ram[15'h1453] =  8'hD7;
		ram[15'h1454] =  8'hFF;
		ram[15'h1455] =  8'h00;
		ram[15'h1456] =  8'h00;
		ram[15'h1457] =  8'hC9;
		ram[15'h1458] =  8'h26;
		ram[15'h1459] =  8'h2D;
		ram[15'h145A] =  8'hE5;
		ram[15'h145B] =  8'h6C;
		ram[15'h145C] =  8'h64;
		ram[15'h145D] =  8'h20;
		ram[15'h145E] =  8'h61;
		ram[15'h145F] =  8'h2C;
		ram[15'h1460] =  8'h28;
		ram[15'h1461] =  8'h6E;
		ram[15'h1462] =  8'h6E;
		ram[15'h1463] =  8'h6E;
		ram[15'h1464] =  8'h6E;
		ram[15'h1465] =  8'h29;
		ram[15'h1466] =  8'h20;
		ram[15'h1467] =  8'h2F;
		ram[15'h1468] =  8'h20;
		ram[15'h1469] =  8'h6C;
		ram[15'h146A] =  8'h64;
		ram[15'h146B] =  8'h20;
		ram[15'h146C] =  8'h28;
		ram[15'h146D] =  8'h6E;
		ram[15'h146E] =  8'h6E;
		ram[15'h146F] =  8'h6E;
		ram[15'h1470] =  8'h6E;
		ram[15'h1471] =  8'h29;
		ram[15'h1472] =  8'h2C;
		ram[15'h1473] =  8'h61;
		ram[15'h1474] =  8'h2E;
		ram[15'h1475] =  8'h2E;
		ram[15'h1476] =  8'h2E;
		ram[15'h1477] =  8'h2E;
		ram[15'h1478] =  8'h2E;
		ram[15'h1479] =  8'h24;
		ram[15'h147A] =  8'hD7;
		ram[15'h147B] =  8'hED;
		ram[15'h147C] =  8'hA8;
		ram[15'h147D] =  8'h00;
		ram[15'h147E] =  8'h00;
		ram[15'h147F] =  8'h52;
		ram[15'h1480] =  8'h98;
		ram[15'h1481] =  8'hFA;
		ram[15'h1482] =  8'h68;
		ram[15'h1483] =  8'hA1;
		ram[15'h1484] =  8'h66;
		ram[15'h1485] =  8'h3D;
		ram[15'h1486] =  8'h00;
		ram[15'h1487] =  8'h3B;
		ram[15'h1488] =  8'h00;
		ram[15'h1489] =  8'h01;
		ram[15'h148A] =  8'h00;
		ram[15'h148B] =  8'hC1;
		ram[15'h148C] =  8'h68;
		ram[15'h148D] =  8'hB7;
		ram[15'h148E] =  8'h20;
		ram[15'h148F] =  8'h00;
		ram[15'h1490] =  8'h10;
		ram[15'h1491] =  8'h00;
		ram[15'h1492] =  8'h00;
		ram[15'h1493] =  8'h00;
		ram[15'h1494] =  8'h00;
		ram[15'h1495] =  8'h00;
		ram[15'h1496] =  8'h00;
		ram[15'h1497] =  8'h00;
		ram[15'h1498] =  8'h00;
		ram[15'h1499] =  8'h00;
		ram[15'h149A] =  8'h00;
		ram[15'h149B] =  8'h00;
		ram[15'h149C] =  8'h00;
		ram[15'h149D] =  8'h00;
		ram[15'h149E] =  8'h00;
		ram[15'h149F] =  8'h00;
		ram[15'h14A0] =  8'h00;
		ram[15'h14A1] =  8'h00;
		ram[15'h14A2] =  8'h00;
		ram[15'h14A3] =  8'h00;
		ram[15'h14A4] =  8'h00;
		ram[15'h14A5] =  8'h00;
		ram[15'h14A6] =  8'h00;
		ram[15'h14A7] =  8'hFF;
		ram[15'h14A8] =  8'hFF;
		ram[15'h14A9] =  8'h00;
		ram[15'h14AA] =  8'h00;
		ram[15'h14AB] =  8'h00;
		ram[15'h14AC] =  8'h00;
		ram[15'h14AD] =  8'h00;
		ram[15'h14AE] =  8'h00;
		ram[15'h14AF] =  8'h00;
		ram[15'h14B0] =  8'h00;
		ram[15'h14B1] =  8'h00;
		ram[15'h14B2] =  8'h00;
		ram[15'h14B3] =  8'hD7;
		ram[15'h14B4] =  8'h00;
		ram[15'h14B5] =  8'h00;
		ram[15'h14B6] =  8'h00;
		ram[15'h14B7] =  8'h94;
		ram[15'h14B8] =  8'hF4;
		ram[15'h14B9] =  8'h27;
		ram[15'h14BA] =  8'h69;
		ram[15'h14BB] =  8'h6C;
		ram[15'h14BC] =  8'h64;
		ram[15'h14BD] =  8'h64;
		ram[15'h14BE] =  8'h3C;
		ram[15'h14BF] =  8'h72;
		ram[15'h14C0] =  8'h3E;
		ram[15'h14C1] =  8'h20;
		ram[15'h14C2] =  8'h28;
		ram[15'h14C3] =  8'h31;
		ram[15'h14C4] =  8'h29;
		ram[15'h14C5] =  8'h2E;
		ram[15'h14C6] =  8'h2E;
		ram[15'h14C7] =  8'h2E;
		ram[15'h14C8] =  8'h2E;
		ram[15'h14C9] =  8'h2E;
		ram[15'h14CA] =  8'h2E;
		ram[15'h14CB] =  8'h2E;
		ram[15'h14CC] =  8'h2E;
		ram[15'h14CD] =  8'h2E;
		ram[15'h14CE] =  8'h2E;
		ram[15'h14CF] =  8'h2E;
		ram[15'h14D0] =  8'h2E;
		ram[15'h14D1] =  8'h2E;
		ram[15'h14D2] =  8'h2E;
		ram[15'h14D3] =  8'h2E;
		ram[15'h14D4] =  8'h2E;
		ram[15'h14D5] =  8'h2E;
		ram[15'h14D6] =  8'h2E;
		ram[15'h14D7] =  8'h2E;
		ram[15'h14D8] =  8'h2E;
		ram[15'h14D9] =  8'h24;
		ram[15'h14DA] =  8'hD7;
		ram[15'h14DB] =  8'hED;
		ram[15'h14DC] =  8'hA8;
		ram[15'h14DD] =  8'h00;
		ram[15'h14DE] =  8'h00;
		ram[15'h14DF] =  8'h2E;
		ram[15'h14E0] =  8'hF1;
		ram[15'h14E1] =  8'h2A;
		ram[15'h14E2] =  8'hEB;
		ram[15'h14E3] =  8'hBA;
		ram[15'h14E4] =  8'hD5;
		ram[15'h14E5] =  8'h3D;
		ram[15'h14E6] =  8'h00;
		ram[15'h14E7] =  8'h3B;
		ram[15'h14E8] =  8'h00;
		ram[15'h14E9] =  8'h02;
		ram[15'h14EA] =  8'h00;
		ram[15'h14EB] =  8'h47;
		ram[15'h14EC] =  8'hFF;
		ram[15'h14ED] =  8'hE4;
		ram[15'h14EE] =  8'hFB;
		ram[15'h14EF] =  8'h00;
		ram[15'h14F0] =  8'h10;
		ram[15'h14F1] =  8'h00;
		ram[15'h14F2] =  8'h00;
		ram[15'h14F3] =  8'h00;
		ram[15'h14F4] =  8'h00;
		ram[15'h14F5] =  8'h00;
		ram[15'h14F6] =  8'h00;
		ram[15'h14F7] =  8'h00;
		ram[15'h14F8] =  8'h00;
		ram[15'h14F9] =  8'h00;
		ram[15'h14FA] =  8'h00;
		ram[15'h14FB] =  8'h00;
		ram[15'h14FC] =  8'h00;
		ram[15'h14FD] =  8'h00;
		ram[15'h14FE] =  8'h00;
		ram[15'h14FF] =  8'h00;
		ram[15'h1500] =  8'h00;
		ram[15'h1501] =  8'h00;
		ram[15'h1502] =  8'h00;
		ram[15'h1503] =  8'h00;
		ram[15'h1504] =  8'h00;
		ram[15'h1505] =  8'h00;
		ram[15'h1506] =  8'h00;
		ram[15'h1507] =  8'hFF;
		ram[15'h1508] =  8'hFF;
		ram[15'h1509] =  8'h00;
		ram[15'h150A] =  8'h00;
		ram[15'h150B] =  8'h00;
		ram[15'h150C] =  8'h00;
		ram[15'h150D] =  8'h00;
		ram[15'h150E] =  8'h00;
		ram[15'h150F] =  8'h00;
		ram[15'h1510] =  8'h00;
		ram[15'h1511] =  8'h00;
		ram[15'h1512] =  8'h00;
		ram[15'h1513] =  8'hD7;
		ram[15'h1514] =  8'h00;
		ram[15'h1515] =  8'h00;
		ram[15'h1516] =  8'h00;
		ram[15'h1517] =  8'h5A;
		ram[15'h1518] =  8'h90;
		ram[15'h1519] =  8'h7E;
		ram[15'h151A] =  8'hD4;
		ram[15'h151B] =  8'h6C;
		ram[15'h151C] =  8'h64;
		ram[15'h151D] =  8'h64;
		ram[15'h151E] =  8'h3C;
		ram[15'h151F] =  8'h72;
		ram[15'h1520] =  8'h3E;
		ram[15'h1521] =  8'h20;
		ram[15'h1522] =  8'h28;
		ram[15'h1523] =  8'h32;
		ram[15'h1524] =  8'h29;
		ram[15'h1525] =  8'h2E;
		ram[15'h1526] =  8'h2E;
		ram[15'h1527] =  8'h2E;
		ram[15'h1528] =  8'h2E;
		ram[15'h1529] =  8'h2E;
		ram[15'h152A] =  8'h2E;
		ram[15'h152B] =  8'h2E;
		ram[15'h152C] =  8'h2E;
		ram[15'h152D] =  8'h2E;
		ram[15'h152E] =  8'h2E;
		ram[15'h152F] =  8'h2E;
		ram[15'h1530] =  8'h2E;
		ram[15'h1531] =  8'h2E;
		ram[15'h1532] =  8'h2E;
		ram[15'h1533] =  8'h2E;
		ram[15'h1534] =  8'h2E;
		ram[15'h1535] =  8'h2E;
		ram[15'h1536] =  8'h2E;
		ram[15'h1537] =  8'h2E;
		ram[15'h1538] =  8'h2E;
		ram[15'h1539] =  8'h24;
		ram[15'h153A] =  8'hD7;
		ram[15'h153B] =  8'hED;
		ram[15'h153C] =  8'hA0;
		ram[15'h153D] =  8'h00;
		ram[15'h153E] =  8'h00;
		ram[15'h153F] =  8'h30;
		ram[15'h1540] =  8'hFE;
		ram[15'h1541] =  8'hCD;
		ram[15'h1542] =  8'h03;
		ram[15'h1543] =  8'h58;
		ram[15'h1544] =  8'h60;
		ram[15'h1545] =  8'h3C;
		ram[15'h1546] =  8'h00;
		ram[15'h1547] =  8'h3A;
		ram[15'h1548] =  8'h00;
		ram[15'h1549] =  8'h01;
		ram[15'h154A] =  8'h00;
		ram[15'h154B] =  8'h04;
		ram[15'h154C] =  8'h60;
		ram[15'h154D] =  8'h88;
		ram[15'h154E] =  8'h26;
		ram[15'h154F] =  8'h00;
		ram[15'h1550] =  8'h10;
		ram[15'h1551] =  8'h00;
		ram[15'h1552] =  8'h00;
		ram[15'h1553] =  8'h00;
		ram[15'h1554] =  8'h00;
		ram[15'h1555] =  8'h00;
		ram[15'h1556] =  8'h00;
		ram[15'h1557] =  8'h00;
		ram[15'h1558] =  8'h00;
		ram[15'h1559] =  8'h00;
		ram[15'h155A] =  8'h00;
		ram[15'h155B] =  8'h00;
		ram[15'h155C] =  8'h00;
		ram[15'h155D] =  8'h00;
		ram[15'h155E] =  8'h00;
		ram[15'h155F] =  8'h00;
		ram[15'h1560] =  8'h00;
		ram[15'h1561] =  8'h00;
		ram[15'h1562] =  8'h00;
		ram[15'h1563] =  8'h00;
		ram[15'h1564] =  8'h00;
		ram[15'h1565] =  8'h00;
		ram[15'h1566] =  8'h00;
		ram[15'h1567] =  8'hFF;
		ram[15'h1568] =  8'hFF;
		ram[15'h1569] =  8'h00;
		ram[15'h156A] =  8'h00;
		ram[15'h156B] =  8'h00;
		ram[15'h156C] =  8'h00;
		ram[15'h156D] =  8'h00;
		ram[15'h156E] =  8'h00;
		ram[15'h156F] =  8'h00;
		ram[15'h1570] =  8'h00;
		ram[15'h1571] =  8'h00;
		ram[15'h1572] =  8'h00;
		ram[15'h1573] =  8'hD7;
		ram[15'h1574] =  8'h00;
		ram[15'h1575] =  8'h00;
		ram[15'h1576] =  8'h00;
		ram[15'h1577] =  8'h9A;
		ram[15'h1578] =  8'hBD;
		ram[15'h1579] =  8'hF6;
		ram[15'h157A] =  8'hB5;
		ram[15'h157B] =  8'h6C;
		ram[15'h157C] =  8'h64;
		ram[15'h157D] =  8'h69;
		ram[15'h157E] =  8'h3C;
		ram[15'h157F] =  8'h72;
		ram[15'h1580] =  8'h3E;
		ram[15'h1581] =  8'h20;
		ram[15'h1582] =  8'h28;
		ram[15'h1583] =  8'h31;
		ram[15'h1584] =  8'h29;
		ram[15'h1585] =  8'h2E;
		ram[15'h1586] =  8'h2E;
		ram[15'h1587] =  8'h2E;
		ram[15'h1588] =  8'h2E;
		ram[15'h1589] =  8'h2E;
		ram[15'h158A] =  8'h2E;
		ram[15'h158B] =  8'h2E;
		ram[15'h158C] =  8'h2E;
		ram[15'h158D] =  8'h2E;
		ram[15'h158E] =  8'h2E;
		ram[15'h158F] =  8'h2E;
		ram[15'h1590] =  8'h2E;
		ram[15'h1591] =  8'h2E;
		ram[15'h1592] =  8'h2E;
		ram[15'h1593] =  8'h2E;
		ram[15'h1594] =  8'h2E;
		ram[15'h1595] =  8'h2E;
		ram[15'h1596] =  8'h2E;
		ram[15'h1597] =  8'h2E;
		ram[15'h1598] =  8'h2E;
		ram[15'h1599] =  8'h24;
		ram[15'h159A] =  8'hD7;
		ram[15'h159B] =  8'hED;
		ram[15'h159C] =  8'hA0;
		ram[15'h159D] =  8'h00;
		ram[15'h159E] =  8'h00;
		ram[15'h159F] =  8'hCE;
		ram[15'h15A0] =  8'h4A;
		ram[15'h15A1] =  8'h6E;
		ram[15'h15A2] =  8'hC2;
		ram[15'h15A3] =  8'h88;
		ram[15'h15A4] =  8'hB1;
		ram[15'h15A5] =  8'h3C;
		ram[15'h15A6] =  8'h00;
		ram[15'h15A7] =  8'h3A;
		ram[15'h15A8] =  8'h00;
		ram[15'h15A9] =  8'h02;
		ram[15'h15AA] =  8'h00;
		ram[15'h15AB] =  8'h14;
		ram[15'h15AC] =  8'h2D;
		ram[15'h15AD] =  8'h9F;
		ram[15'h15AE] =  8'hA3;
		ram[15'h15AF] =  8'h00;
		ram[15'h15B0] =  8'h10;
		ram[15'h15B1] =  8'h00;
		ram[15'h15B2] =  8'h00;
		ram[15'h15B3] =  8'h00;
		ram[15'h15B4] =  8'h00;
		ram[15'h15B5] =  8'h00;
		ram[15'h15B6] =  8'h00;
		ram[15'h15B7] =  8'h00;
		ram[15'h15B8] =  8'h00;
		ram[15'h15B9] =  8'h00;
		ram[15'h15BA] =  8'h00;
		ram[15'h15BB] =  8'h00;
		ram[15'h15BC] =  8'h00;
		ram[15'h15BD] =  8'h00;
		ram[15'h15BE] =  8'h00;
		ram[15'h15BF] =  8'h00;
		ram[15'h15C0] =  8'h00;
		ram[15'h15C1] =  8'h00;
		ram[15'h15C2] =  8'h00;
		ram[15'h15C3] =  8'h00;
		ram[15'h15C4] =  8'h00;
		ram[15'h15C5] =  8'h00;
		ram[15'h15C6] =  8'h00;
		ram[15'h15C7] =  8'hFF;
		ram[15'h15C8] =  8'hFF;
		ram[15'h15C9] =  8'h00;
		ram[15'h15CA] =  8'h00;
		ram[15'h15CB] =  8'h00;
		ram[15'h15CC] =  8'h00;
		ram[15'h15CD] =  8'h00;
		ram[15'h15CE] =  8'h00;
		ram[15'h15CF] =  8'h00;
		ram[15'h15D0] =  8'h00;
		ram[15'h15D1] =  8'h00;
		ram[15'h15D2] =  8'h00;
		ram[15'h15D3] =  8'hD7;
		ram[15'h15D4] =  8'h00;
		ram[15'h15D5] =  8'h00;
		ram[15'h15D6] =  8'h00;
		ram[15'h15D7] =  8'hEB;
		ram[15'h15D8] =  8'h59;
		ram[15'h15D9] =  8'h89;
		ram[15'h15DA] =  8'h1B;
		ram[15'h15DB] =  8'h6C;
		ram[15'h15DC] =  8'h64;
		ram[15'h15DD] =  8'h69;
		ram[15'h15DE] =  8'h3C;
		ram[15'h15DF] =  8'h72;
		ram[15'h15E0] =  8'h3E;
		ram[15'h15E1] =  8'h20;
		ram[15'h15E2] =  8'h28;
		ram[15'h15E3] =  8'h32;
		ram[15'h15E4] =  8'h29;
		ram[15'h15E5] =  8'h2E;
		ram[15'h15E6] =  8'h2E;
		ram[15'h15E7] =  8'h2E;
		ram[15'h15E8] =  8'h2E;
		ram[15'h15E9] =  8'h2E;
		ram[15'h15EA] =  8'h2E;
		ram[15'h15EB] =  8'h2E;
		ram[15'h15EC] =  8'h2E;
		ram[15'h15ED] =  8'h2E;
		ram[15'h15EE] =  8'h2E;
		ram[15'h15EF] =  8'h2E;
		ram[15'h15F0] =  8'h2E;
		ram[15'h15F1] =  8'h2E;
		ram[15'h15F2] =  8'h2E;
		ram[15'h15F3] =  8'h2E;
		ram[15'h15F4] =  8'h2E;
		ram[15'h15F5] =  8'h2E;
		ram[15'h15F6] =  8'h2E;
		ram[15'h15F7] =  8'h2E;
		ram[15'h15F8] =  8'h2E;
		ram[15'h15F9] =  8'h24;
		ram[15'h15FA] =  8'hD7;
		ram[15'h15FB] =  8'hED;
		ram[15'h15FC] =  8'h44;
		ram[15'h15FD] =  8'h00;
		ram[15'h15FE] =  8'h00;
		ram[15'h15FF] =  8'hA2;
		ram[15'h1600] =  8'h38;
		ram[15'h1601] =  8'h6B;
		ram[15'h1602] =  8'h5F;
		ram[15'h1603] =  8'h34;
		ram[15'h1604] =  8'hD9;
		ram[15'h1605] =  8'hE4;
		ram[15'h1606] =  8'h57;
		ram[15'h1607] =  8'hD6;
		ram[15'h1608] =  8'hD2;
		ram[15'h1609] =  8'h42;
		ram[15'h160A] =  8'h46;
		ram[15'h160B] =  8'h43;
		ram[15'h160C] =  8'h5A;
		ram[15'h160D] =  8'hCC;
		ram[15'h160E] =  8'h09;
		ram[15'h160F] =  8'h00;
		ram[15'h1610] =  8'h00;
		ram[15'h1611] =  8'h00;
		ram[15'h1612] =  8'h00;
		ram[15'h1613] =  8'h00;
		ram[15'h1614] =  8'h00;
		ram[15'h1615] =  8'h00;
		ram[15'h1616] =  8'h00;
		ram[15'h1617] =  8'h00;
		ram[15'h1618] =  8'h00;
		ram[15'h1619] =  8'h00;
		ram[15'h161A] =  8'h00;
		ram[15'h161B] =  8'h00;
		ram[15'h161C] =  8'h00;
		ram[15'h161D] =  8'h00;
		ram[15'h161E] =  8'h00;
		ram[15'h161F] =  8'hD7;
		ram[15'h1620] =  8'hFF;
		ram[15'h1621] =  8'h00;
		ram[15'h1622] =  8'h00;
		ram[15'h1623] =  8'h00;
		ram[15'h1624] =  8'h00;
		ram[15'h1625] =  8'h00;
		ram[15'h1626] =  8'h00;
		ram[15'h1627] =  8'h00;
		ram[15'h1628] =  8'h00;
		ram[15'h1629] =  8'h00;
		ram[15'h162A] =  8'h00;
		ram[15'h162B] =  8'h00;
		ram[15'h162C] =  8'h00;
		ram[15'h162D] =  8'h00;
		ram[15'h162E] =  8'h00;
		ram[15'h162F] =  8'h00;
		ram[15'h1630] =  8'h00;
		ram[15'h1631] =  8'h00;
		ram[15'h1632] =  8'h00;
		ram[15'h1633] =  8'h00;
		ram[15'h1634] =  8'h00;
		ram[15'h1635] =  8'h00;
		ram[15'h1636] =  8'h00;
		ram[15'h1637] =  8'h6A;
		ram[15'h1638] =  8'h3C;
		ram[15'h1639] =  8'h3B;
		ram[15'h163A] =  8'hBD;
		ram[15'h163B] =  8'h6E;
		ram[15'h163C] =  8'h65;
		ram[15'h163D] =  8'h67;
		ram[15'h163E] =  8'h2E;
		ram[15'h163F] =  8'h2E;
		ram[15'h1640] =  8'h2E;
		ram[15'h1641] =  8'h2E;
		ram[15'h1642] =  8'h2E;
		ram[15'h1643] =  8'h2E;
		ram[15'h1644] =  8'h2E;
		ram[15'h1645] =  8'h2E;
		ram[15'h1646] =  8'h2E;
		ram[15'h1647] =  8'h2E;
		ram[15'h1648] =  8'h2E;
		ram[15'h1649] =  8'h2E;
		ram[15'h164A] =  8'h2E;
		ram[15'h164B] =  8'h2E;
		ram[15'h164C] =  8'h2E;
		ram[15'h164D] =  8'h2E;
		ram[15'h164E] =  8'h2E;
		ram[15'h164F] =  8'h2E;
		ram[15'h1650] =  8'h2E;
		ram[15'h1651] =  8'h2E;
		ram[15'h1652] =  8'h2E;
		ram[15'h1653] =  8'h2E;
		ram[15'h1654] =  8'h2E;
		ram[15'h1655] =  8'h2E;
		ram[15'h1656] =  8'h2E;
		ram[15'h1657] =  8'h2E;
		ram[15'h1658] =  8'h2E;
		ram[15'h1659] =  8'h24;
		ram[15'h165A] =  8'hD7;
		ram[15'h165B] =  8'hED;
		ram[15'h165C] =  8'h67;
		ram[15'h165D] =  8'h00;
		ram[15'h165E] =  8'h00;
		ram[15'h165F] =  8'hCB;
		ram[15'h1660] =  8'h91;
		ram[15'h1661] =  8'h8B;
		ram[15'h1662] =  8'hC4;
		ram[15'h1663] =  8'h62;
		ram[15'h1664] =  8'hFA;
		ram[15'h1665] =  8'h3A;
		ram[15'h1666] =  8'h00;
		ram[15'h1667] =  8'h20;
		ram[15'h1668] =  8'hE7;
		ram[15'h1669] =  8'h79;
		ram[15'h166A] =  8'hB4;
		ram[15'h166B] =  8'h40;
		ram[15'h166C] =  8'h06;
		ram[15'h166D] =  8'hE2;
		ram[15'h166E] =  8'h8A;
		ram[15'h166F] =  8'h00;
		ram[15'h1670] =  8'h08;
		ram[15'h1671] =  8'h00;
		ram[15'h1672] =  8'h00;
		ram[15'h1673] =  8'hFF;
		ram[15'h1674] =  8'h00;
		ram[15'h1675] =  8'h00;
		ram[15'h1676] =  8'h00;
		ram[15'h1677] =  8'h00;
		ram[15'h1678] =  8'h00;
		ram[15'h1679] =  8'h00;
		ram[15'h167A] =  8'h00;
		ram[15'h167B] =  8'h00;
		ram[15'h167C] =  8'h00;
		ram[15'h167D] =  8'h00;
		ram[15'h167E] =  8'h00;
		ram[15'h167F] =  8'h00;
		ram[15'h1680] =  8'h00;
		ram[15'h1681] =  8'h00;
		ram[15'h1682] =  8'h00;
		ram[15'h1683] =  8'h00;
		ram[15'h1684] =  8'h00;
		ram[15'h1685] =  8'h00;
		ram[15'h1686] =  8'h00;
		ram[15'h1687] =  8'h00;
		ram[15'h1688] =  8'h00;
		ram[15'h1689] =  8'h00;
		ram[15'h168A] =  8'h00;
		ram[15'h168B] =  8'h00;
		ram[15'h168C] =  8'h00;
		ram[15'h168D] =  8'h00;
		ram[15'h168E] =  8'h00;
		ram[15'h168F] =  8'h00;
		ram[15'h1690] =  8'h00;
		ram[15'h1691] =  8'h00;
		ram[15'h1692] =  8'h00;
		ram[15'h1693] =  8'hD7;
		ram[15'h1694] =  8'hFF;
		ram[15'h1695] =  8'h00;
		ram[15'h1696] =  8'h00;
		ram[15'h1697] =  8'h95;
		ram[15'h1698] =  8'h5B;
		ram[15'h1699] =  8'hA3;
		ram[15'h169A] =  8'h26;
		ram[15'h169B] =  8'h3C;
		ram[15'h169C] =  8'h72;
		ram[15'h169D] =  8'h72;
		ram[15'h169E] =  8'h64;
		ram[15'h169F] =  8'h2C;
		ram[15'h16A0] =  8'h72;
		ram[15'h16A1] =  8'h6C;
		ram[15'h16A2] =  8'h64;
		ram[15'h16A3] =  8'h3E;
		ram[15'h16A4] =  8'h2E;
		ram[15'h16A5] =  8'h2E;
		ram[15'h16A6] =  8'h2E;
		ram[15'h16A7] =  8'h2E;
		ram[15'h16A8] =  8'h2E;
		ram[15'h16A9] =  8'h2E;
		ram[15'h16AA] =  8'h2E;
		ram[15'h16AB] =  8'h2E;
		ram[15'h16AC] =  8'h2E;
		ram[15'h16AD] =  8'h2E;
		ram[15'h16AE] =  8'h2E;
		ram[15'h16AF] =  8'h2E;
		ram[15'h16B0] =  8'h2E;
		ram[15'h16B1] =  8'h2E;
		ram[15'h16B2] =  8'h2E;
		ram[15'h16B3] =  8'h2E;
		ram[15'h16B4] =  8'h2E;
		ram[15'h16B5] =  8'h2E;
		ram[15'h16B6] =  8'h2E;
		ram[15'h16B7] =  8'h2E;
		ram[15'h16B8] =  8'h2E;
		ram[15'h16B9] =  8'h24;
		ram[15'h16BA] =  8'hD7;
		ram[15'h16BB] =  8'h07;
		ram[15'h16BC] =  8'h00;
		ram[15'h16BD] =  8'h00;
		ram[15'h16BE] =  8'h00;
		ram[15'h16BF] =  8'h92;
		ram[15'h16C0] =  8'hCB;
		ram[15'h16C1] =  8'h43;
		ram[15'h16C2] =  8'h6D;
		ram[15'h16C3] =  8'h90;
		ram[15'h16C4] =  8'h0A;
		ram[15'h16C5] =  8'h84;
		ram[15'h16C6] =  8'hC2;
		ram[15'h16C7] =  8'h53;
		ram[15'h16C8] =  8'h0C;
		ram[15'h16C9] =  8'h0E;
		ram[15'h16CA] =  8'hF5;
		ram[15'h16CB] =  8'h91;
		ram[15'h16CC] =  8'hEB;
		ram[15'h16CD] =  8'hFC;
		ram[15'h16CE] =  8'h40;
		ram[15'h16CF] =  8'h18;
		ram[15'h16D0] =  8'h00;
		ram[15'h16D1] =  8'h00;
		ram[15'h16D2] =  8'h00;
		ram[15'h16D3] =  8'h00;
		ram[15'h16D4] =  8'h00;
		ram[15'h16D5] =  8'h00;
		ram[15'h16D6] =  8'h00;
		ram[15'h16D7] =  8'h00;
		ram[15'h16D8] =  8'h00;
		ram[15'h16D9] =  8'h00;
		ram[15'h16DA] =  8'h00;
		ram[15'h16DB] =  8'h00;
		ram[15'h16DC] =  8'h00;
		ram[15'h16DD] =  8'h00;
		ram[15'h16DE] =  8'h00;
		ram[15'h16DF] =  8'h00;
		ram[15'h16E0] =  8'hFF;
		ram[15'h16E1] =  8'h00;
		ram[15'h16E2] =  8'h00;
		ram[15'h16E3] =  8'h00;
		ram[15'h16E4] =  8'h00;
		ram[15'h16E5] =  8'h00;
		ram[15'h16E6] =  8'h00;
		ram[15'h16E7] =  8'h00;
		ram[15'h16E8] =  8'h00;
		ram[15'h16E9] =  8'h00;
		ram[15'h16EA] =  8'h00;
		ram[15'h16EB] =  8'h00;
		ram[15'h16EC] =  8'h00;
		ram[15'h16ED] =  8'h00;
		ram[15'h16EE] =  8'h00;
		ram[15'h16EF] =  8'h00;
		ram[15'h16F0] =  8'h00;
		ram[15'h16F1] =  8'h00;
		ram[15'h16F2] =  8'h00;
		ram[15'h16F3] =  8'hD7;
		ram[15'h16F4] =  8'h00;
		ram[15'h16F5] =  8'h00;
		ram[15'h16F6] =  8'h00;
		ram[15'h16F7] =  8'h25;
		ram[15'h16F8] =  8'h13;
		ram[15'h16F9] =  8'h30;
		ram[15'h16FA] =  8'hAE;
		ram[15'h16FB] =  8'h3C;
		ram[15'h16FC] =  8'h72;
		ram[15'h16FD] =  8'h6C;
		ram[15'h16FE] =  8'h63;
		ram[15'h16FF] =  8'h61;
		ram[15'h1700] =  8'h2C;
		ram[15'h1701] =  8'h72;
		ram[15'h1702] =  8'h72;
		ram[15'h1703] =  8'h63;
		ram[15'h1704] =  8'h61;
		ram[15'h1705] =  8'h2C;
		ram[15'h1706] =  8'h72;
		ram[15'h1707] =  8'h6C;
		ram[15'h1708] =  8'h61;
		ram[15'h1709] =  8'h2C;
		ram[15'h170A] =  8'h72;
		ram[15'h170B] =  8'h72;
		ram[15'h170C] =  8'h61;
		ram[15'h170D] =  8'h3E;
		ram[15'h170E] =  8'h2E;
		ram[15'h170F] =  8'h2E;
		ram[15'h1710] =  8'h2E;
		ram[15'h1711] =  8'h2E;
		ram[15'h1712] =  8'h2E;
		ram[15'h1713] =  8'h2E;
		ram[15'h1714] =  8'h2E;
		ram[15'h1715] =  8'h2E;
		ram[15'h1716] =  8'h2E;
		ram[15'h1717] =  8'h2E;
		ram[15'h1718] =  8'h2E;
		ram[15'h1719] =  8'h24;
		ram[15'h171A] =  8'hD7;
		ram[15'h171B] =  8'hDD;
		ram[15'h171C] =  8'hCB;
		ram[15'h171D] =  8'h01;
		ram[15'h171E] =  8'h06;
		ram[15'h171F] =  8'hAF;
		ram[15'h1720] =  8'hDD;
		ram[15'h1721] =  8'h39;
		ram[15'h1722] =  8'h00;
		ram[15'h1723] =  8'h39;
		ram[15'h1724] =  8'h00;
		ram[15'h1725] =  8'h3C;
		ram[15'h1726] =  8'hFF;
		ram[15'h1727] =  8'hF6;
		ram[15'h1728] =  8'hDB;
		ram[15'h1729] =  8'hF4;
		ram[15'h172A] =  8'h94;
		ram[15'h172B] =  8'h82;
		ram[15'h172C] =  8'h80;
		ram[15'h172D] =  8'hD9;
		ram[15'h172E] =  8'h61;
		ram[15'h172F] =  8'h20;
		ram[15'h1730] =  8'h00;
		ram[15'h1731] =  8'h00;
		ram[15'h1732] =  8'h38;
		ram[15'h1733] =  8'h00;
		ram[15'h1734] =  8'h00;
		ram[15'h1735] =  8'h00;
		ram[15'h1736] =  8'h00;
		ram[15'h1737] =  8'h00;
		ram[15'h1738] =  8'h00;
		ram[15'h1739] =  8'h00;
		ram[15'h173A] =  8'h00;
		ram[15'h173B] =  8'h00;
		ram[15'h173C] =  8'h00;
		ram[15'h173D] =  8'h00;
		ram[15'h173E] =  8'h00;
		ram[15'h173F] =  8'h80;
		ram[15'h1740] =  8'h00;
		ram[15'h1741] =  8'h00;
		ram[15'h1742] =  8'h00;
		ram[15'h1743] =  8'h00;
		ram[15'h1744] =  8'h00;
		ram[15'h1745] =  8'h00;
		ram[15'h1746] =  8'h00;
		ram[15'h1747] =  8'hFF;
		ram[15'h1748] =  8'h00;
		ram[15'h1749] =  8'h00;
		ram[15'h174A] =  8'h00;
		ram[15'h174B] =  8'h00;
		ram[15'h174C] =  8'h00;
		ram[15'h174D] =  8'h00;
		ram[15'h174E] =  8'h00;
		ram[15'h174F] =  8'h00;
		ram[15'h1750] =  8'h00;
		ram[15'h1751] =  8'h00;
		ram[15'h1752] =  8'h00;
		ram[15'h1753] =  8'h57;
		ram[15'h1754] =  8'h00;
		ram[15'h1755] =  8'h00;
		ram[15'h1756] =  8'h00;
		ram[15'h1757] =  8'h71;
		ram[15'h1758] =  8'h3A;
		ram[15'h1759] =  8'hCD;
		ram[15'h175A] =  8'h81;
		ram[15'h175B] =  8'h73;
		ram[15'h175C] =  8'h68;
		ram[15'h175D] =  8'h66;
		ram[15'h175E] =  8'h2F;
		ram[15'h175F] =  8'h72;
		ram[15'h1760] =  8'h6F;
		ram[15'h1761] =  8'h74;
		ram[15'h1762] =  8'h20;
		ram[15'h1763] =  8'h28;
		ram[15'h1764] =  8'h3C;
		ram[15'h1765] =  8'h69;
		ram[15'h1766] =  8'h78;
		ram[15'h1767] =  8'h2C;
		ram[15'h1768] =  8'h69;
		ram[15'h1769] =  8'h79;
		ram[15'h176A] =  8'h3E;
		ram[15'h176B] =  8'h2B;
		ram[15'h176C] =  8'h31;
		ram[15'h176D] =  8'h29;
		ram[15'h176E] =  8'h2E;
		ram[15'h176F] =  8'h2E;
		ram[15'h1770] =  8'h2E;
		ram[15'h1771] =  8'h2E;
		ram[15'h1772] =  8'h2E;
		ram[15'h1773] =  8'h2E;
		ram[15'h1774] =  8'h2E;
		ram[15'h1775] =  8'h2E;
		ram[15'h1776] =  8'h2E;
		ram[15'h1777] =  8'h2E;
		ram[15'h1778] =  8'h2E;
		ram[15'h1779] =  8'h24;
		ram[15'h177A] =  8'hD7;
		ram[15'h177B] =  8'hCB;
		ram[15'h177C] =  8'h00;
		ram[15'h177D] =  8'h00;
		ram[15'h177E] =  8'h00;
		ram[15'h177F] =  8'hEB;
		ram[15'h1780] =  8'hCC;
		ram[15'h1781] =  8'h4A;
		ram[15'h1782] =  8'h5D;
		ram[15'h1783] =  8'h07;
		ram[15'h1784] =  8'hE0;
		ram[15'h1785] =  8'h3A;
		ram[15'h1786] =  8'h00;
		ram[15'h1787] =  8'h95;
		ram[15'h1788] =  8'h13;
		ram[15'h1789] =  8'hEE;
		ram[15'h178A] =  8'h30;
		ram[15'h178B] =  8'h43;
		ram[15'h178C] =  8'h78;
		ram[15'h178D] =  8'hAD;
		ram[15'h178E] =  8'h3D;
		ram[15'h178F] =  8'h00;
		ram[15'h1790] =  8'h3F;
		ram[15'h1791] =  8'h00;
		ram[15'h1792] =  8'h00;
		ram[15'h1793] =  8'h00;
		ram[15'h1794] =  8'h00;
		ram[15'h1795] =  8'h00;
		ram[15'h1796] =  8'h00;
		ram[15'h1797] =  8'h00;
		ram[15'h1798] =  8'h00;
		ram[15'h1799] =  8'h00;
		ram[15'h179A] =  8'h00;
		ram[15'h179B] =  8'h00;
		ram[15'h179C] =  8'h00;
		ram[15'h179D] =  8'h00;
		ram[15'h179E] =  8'h00;
		ram[15'h179F] =  8'h80;
		ram[15'h17A0] =  8'h00;
		ram[15'h17A1] =  8'h00;
		ram[15'h17A2] =  8'h00;
		ram[15'h17A3] =  8'h00;
		ram[15'h17A4] =  8'h00;
		ram[15'h17A5] =  8'h00;
		ram[15'h17A6] =  8'h00;
		ram[15'h17A7] =  8'hFF;
		ram[15'h17A8] =  8'h00;
		ram[15'h17A9] =  8'h00;
		ram[15'h17AA] =  8'h00;
		ram[15'h17AB] =  8'h00;
		ram[15'h17AC] =  8'h00;
		ram[15'h17AD] =  8'h00;
		ram[15'h17AE] =  8'h00;
		ram[15'h17AF] =  8'hFF;
		ram[15'h17B0] =  8'hFF;
		ram[15'h17B1] =  8'hFF;
		ram[15'h17B2] =  8'hFF;
		ram[15'h17B3] =  8'h57;
		ram[15'h17B4] =  8'hFF;
		ram[15'h17B5] =  8'h00;
		ram[15'h17B6] =  8'h00;
		ram[15'h17B7] =  8'hEB;
		ram[15'h17B8] =  8'h60;
		ram[15'h17B9] =  8'h4D;
		ram[15'h17BA] =  8'h58;
		ram[15'h17BB] =  8'h73;
		ram[15'h17BC] =  8'h68;
		ram[15'h17BD] =  8'h66;
		ram[15'h17BE] =  8'h2F;
		ram[15'h17BF] =  8'h72;
		ram[15'h17C0] =  8'h6F;
		ram[15'h17C1] =  8'h74;
		ram[15'h17C2] =  8'h20;
		ram[15'h17C3] =  8'h3C;
		ram[15'h17C4] =  8'h62;
		ram[15'h17C5] =  8'h2C;
		ram[15'h17C6] =  8'h63;
		ram[15'h17C7] =  8'h2C;
		ram[15'h17C8] =  8'h64;
		ram[15'h17C9] =  8'h2C;
		ram[15'h17CA] =  8'h65;
		ram[15'h17CB] =  8'h2C;
		ram[15'h17CC] =  8'h68;
		ram[15'h17CD] =  8'h2C;
		ram[15'h17CE] =  8'h6C;
		ram[15'h17CF] =  8'h2C;
		ram[15'h17D0] =  8'h28;
		ram[15'h17D1] =  8'h68;
		ram[15'h17D2] =  8'h6C;
		ram[15'h17D3] =  8'h29;
		ram[15'h17D4] =  8'h2C;
		ram[15'h17D5] =  8'h61;
		ram[15'h17D6] =  8'h3E;
		ram[15'h17D7] =  8'h2E;
		ram[15'h17D8] =  8'h2E;
		ram[15'h17D9] =  8'h24;
		ram[15'h17DA] =  8'hD7;
		ram[15'h17DB] =  8'hCB;
		ram[15'h17DC] =  8'h80;
		ram[15'h17DD] =  8'h00;
		ram[15'h17DE] =  8'h00;
		ram[15'h17DF] =  8'hD5;
		ram[15'h17E0] =  8'h2C;
		ram[15'h17E1] =  8'hAB;
		ram[15'h17E2] =  8'h97;
		ram[15'h17E3] =  8'hFF;
		ram[15'h17E4] =  8'h39;
		ram[15'h17E5] =  8'h3A;
		ram[15'h17E6] =  8'h00;
		ram[15'h17E7] =  8'h4B;
		ram[15'h17E8] =  8'hD1;
		ram[15'h17E9] =  8'hB2;
		ram[15'h17EA] =  8'h6A;
		ram[15'h17EB] =  8'h53;
		ram[15'h17EC] =  8'h27;
		ram[15'h17ED] =  8'h38;
		ram[15'h17EE] =  8'hB5;
		ram[15'h17EF] =  8'h00;
		ram[15'h17F0] =  8'h7F;
		ram[15'h17F1] =  8'h00;
		ram[15'h17F2] =  8'h00;
		ram[15'h17F3] =  8'h00;
		ram[15'h17F4] =  8'h00;
		ram[15'h17F5] =  8'h00;
		ram[15'h17F6] =  8'h00;
		ram[15'h17F7] =  8'h00;
		ram[15'h17F8] =  8'h00;
		ram[15'h17F9] =  8'h00;
		ram[15'h17FA] =  8'h00;
		ram[15'h17FB] =  8'h00;
		ram[15'h17FC] =  8'h00;
		ram[15'h17FD] =  8'h00;
		ram[15'h17FE] =  8'h00;
		ram[15'h17FF] =  8'h00;
		ram[15'h1800] =  8'h00;
		ram[15'h1801] =  8'h00;
		ram[15'h1802] =  8'h00;
		ram[15'h1803] =  8'h00;
		ram[15'h1804] =  8'h00;
		ram[15'h1805] =  8'h00;
		ram[15'h1806] =  8'h00;
		ram[15'h1807] =  8'hFF;
		ram[15'h1808] =  8'h00;
		ram[15'h1809] =  8'h00;
		ram[15'h180A] =  8'h00;
		ram[15'h180B] =  8'h00;
		ram[15'h180C] =  8'h00;
		ram[15'h180D] =  8'h00;
		ram[15'h180E] =  8'h00;
		ram[15'h180F] =  8'hFF;
		ram[15'h1810] =  8'hFF;
		ram[15'h1811] =  8'hFF;
		ram[15'h1812] =  8'hFF;
		ram[15'h1813] =  8'hD7;
		ram[15'h1814] =  8'hFF;
		ram[15'h1815] =  8'h00;
		ram[15'h1816] =  8'h00;
		ram[15'h1817] =  8'h8B;
		ram[15'h1818] =  8'h57;
		ram[15'h1819] =  8'hF0;
		ram[15'h181A] =  8'h08;
		ram[15'h181B] =  8'h3C;
		ram[15'h181C] =  8'h73;
		ram[15'h181D] =  8'h65;
		ram[15'h181E] =  8'h74;
		ram[15'h181F] =  8'h2C;
		ram[15'h1820] =  8'h72;
		ram[15'h1821] =  8'h65;
		ram[15'h1822] =  8'h73;
		ram[15'h1823] =  8'h3E;
		ram[15'h1824] =  8'h20;
		ram[15'h1825] =  8'h6E;
		ram[15'h1826] =  8'h2C;
		ram[15'h1827] =  8'h3C;
		ram[15'h1828] =  8'h62;
		ram[15'h1829] =  8'h63;
		ram[15'h182A] =  8'h64;
		ram[15'h182B] =  8'h65;
		ram[15'h182C] =  8'h68;
		ram[15'h182D] =  8'h6C;
		ram[15'h182E] =  8'h28;
		ram[15'h182F] =  8'h68;
		ram[15'h1830] =  8'h6C;
		ram[15'h1831] =  8'h29;
		ram[15'h1832] =  8'h61;
		ram[15'h1833] =  8'h3E;
		ram[15'h1834] =  8'h2E;
		ram[15'h1835] =  8'h2E;
		ram[15'h1836] =  8'h2E;
		ram[15'h1837] =  8'h2E;
		ram[15'h1838] =  8'h2E;
		ram[15'h1839] =  8'h24;
		ram[15'h183A] =  8'hD7;
		ram[15'h183B] =  8'hDD;
		ram[15'h183C] =  8'hCB;
		ram[15'h183D] =  8'h01;
		ram[15'h183E] =  8'h86;
		ram[15'h183F] =  8'h44;
		ram[15'h1840] =  8'hFB;
		ram[15'h1841] =  8'h39;
		ram[15'h1842] =  8'h00;
		ram[15'h1843] =  8'h39;
		ram[15'h1844] =  8'h00;
		ram[15'h1845] =  8'h09;
		ram[15'h1846] =  8'hBA;
		ram[15'h1847] =  8'hBE;
		ram[15'h1848] =  8'h68;
		ram[15'h1849] =  8'hD8;
		ram[15'h184A] =  8'h32;
		ram[15'h184B] =  8'h10;
		ram[15'h184C] =  8'h5E;
		ram[15'h184D] =  8'h67;
		ram[15'h184E] =  8'hA8;
		ram[15'h184F] =  8'h20;
		ram[15'h1850] =  8'h00;
		ram[15'h1851] =  8'h00;
		ram[15'h1852] =  8'h78;
		ram[15'h1853] =  8'h00;
		ram[15'h1854] =  8'h00;
		ram[15'h1855] =  8'h00;
		ram[15'h1856] =  8'h00;
		ram[15'h1857] =  8'h00;
		ram[15'h1858] =  8'h00;
		ram[15'h1859] =  8'h00;
		ram[15'h185A] =  8'h00;
		ram[15'h185B] =  8'h00;
		ram[15'h185C] =  8'h00;
		ram[15'h185D] =  8'h00;
		ram[15'h185E] =  8'h00;
		ram[15'h185F] =  8'h00;
		ram[15'h1860] =  8'h00;
		ram[15'h1861] =  8'h00;
		ram[15'h1862] =  8'h00;
		ram[15'h1863] =  8'h00;
		ram[15'h1864] =  8'h00;
		ram[15'h1865] =  8'h00;
		ram[15'h1866] =  8'h00;
		ram[15'h1867] =  8'hFF;
		ram[15'h1868] =  8'h00;
		ram[15'h1869] =  8'h00;
		ram[15'h186A] =  8'h00;
		ram[15'h186B] =  8'h00;
		ram[15'h186C] =  8'h00;
		ram[15'h186D] =  8'h00;
		ram[15'h186E] =  8'h00;
		ram[15'h186F] =  8'h00;
		ram[15'h1870] =  8'h00;
		ram[15'h1871] =  8'h00;
		ram[15'h1872] =  8'h00;
		ram[15'h1873] =  8'hD7;
		ram[15'h1874] =  8'h00;
		ram[15'h1875] =  8'h00;
		ram[15'h1876] =  8'h00;
		ram[15'h1877] =  8'hCC;
		ram[15'h1878] =  8'h63;
		ram[15'h1879] =  8'hF9;
		ram[15'h187A] =  8'h8A;
		ram[15'h187B] =  8'h3C;
		ram[15'h187C] =  8'h73;
		ram[15'h187D] =  8'h65;
		ram[15'h187E] =  8'h74;
		ram[15'h187F] =  8'h2C;
		ram[15'h1880] =  8'h72;
		ram[15'h1881] =  8'h65;
		ram[15'h1882] =  8'h73;
		ram[15'h1883] =  8'h3E;
		ram[15'h1884] =  8'h20;
		ram[15'h1885] =  8'h6E;
		ram[15'h1886] =  8'h2C;
		ram[15'h1887] =  8'h28;
		ram[15'h1888] =  8'h3C;
		ram[15'h1889] =  8'h69;
		ram[15'h188A] =  8'h78;
		ram[15'h188B] =  8'h2C;
		ram[15'h188C] =  8'h69;
		ram[15'h188D] =  8'h79;
		ram[15'h188E] =  8'h3E;
		ram[15'h188F] =  8'h2B;
		ram[15'h1890] =  8'h31;
		ram[15'h1891] =  8'h29;
		ram[15'h1892] =  8'h2E;
		ram[15'h1893] =  8'h2E;
		ram[15'h1894] =  8'h2E;
		ram[15'h1895] =  8'h2E;
		ram[15'h1896] =  8'h2E;
		ram[15'h1897] =  8'h2E;
		ram[15'h1898] =  8'h2E;
		ram[15'h1899] =  8'h24;
		ram[15'h189A] =  8'hD7;
		ram[15'h189B] =  8'hDD;
		ram[15'h189C] =  8'h70;
		ram[15'h189D] =  8'h01;
		ram[15'h189E] =  8'h00;
		ram[15'h189F] =  8'h0D;
		ram[15'h18A0] =  8'h27;
		ram[15'h18A1] =  8'h39;
		ram[15'h18A2] =  8'h00;
		ram[15'h18A3] =  8'h39;
		ram[15'h18A4] =  8'h00;
		ram[15'h18A5] =  8'h3A;
		ram[15'h18A6] =  8'hB7;
		ram[15'h18A7] =  8'h7B;
		ram[15'h18A8] =  8'h88;
		ram[15'h18A9] =  8'hEE;
		ram[15'h18AA] =  8'h99;
		ram[15'h18AB] =  8'h86;
		ram[15'h18AC] =  8'h70;
		ram[15'h18AD] =  8'h07;
		ram[15'h18AE] =  8'hCA;
		ram[15'h18AF] =  8'h20;
		ram[15'h18B0] =  8'h03;
		ram[15'h18B1] =  8'h00;
		ram[15'h18B2] =  8'h00;
		ram[15'h18B3] =  8'h00;
		ram[15'h18B4] =  8'h00;
		ram[15'h18B5] =  8'h01;
		ram[15'h18B6] =  8'h00;
		ram[15'h18B7] =  8'h01;
		ram[15'h18B8] =  8'h00;
		ram[15'h18B9] =  8'h00;
		ram[15'h18BA] =  8'h00;
		ram[15'h18BB] =  8'h00;
		ram[15'h18BC] =  8'h00;
		ram[15'h18BD] =  8'h00;
		ram[15'h18BE] =  8'h00;
		ram[15'h18BF] =  8'h00;
		ram[15'h18C0] =  8'h00;
		ram[15'h18C1] =  8'h00;
		ram[15'h18C2] =  8'h00;
		ram[15'h18C3] =  8'h00;
		ram[15'h18C4] =  8'h00;
		ram[15'h18C5] =  8'h00;
		ram[15'h18C6] =  8'h00;
		ram[15'h18C7] =  8'h00;
		ram[15'h18C8] =  8'h00;
		ram[15'h18C9] =  8'h00;
		ram[15'h18CA] =  8'h00;
		ram[15'h18CB] =  8'h00;
		ram[15'h18CC] =  8'h00;
		ram[15'h18CD] =  8'h00;
		ram[15'h18CE] =  8'h00;
		ram[15'h18CF] =  8'hFF;
		ram[15'h18D0] =  8'hFF;
		ram[15'h18D1] =  8'hFF;
		ram[15'h18D2] =  8'hFF;
		ram[15'h18D3] =  8'h00;
		ram[15'h18D4] =  8'h00;
		ram[15'h18D5] =  8'h00;
		ram[15'h18D6] =  8'h00;
		ram[15'h18D7] =  8'h04;
		ram[15'h18D8] =  8'h62;
		ram[15'h18D9] =  8'h6A;
		ram[15'h18DA] =  8'hBF;
		ram[15'h18DB] =  8'h6C;
		ram[15'h18DC] =  8'h64;
		ram[15'h18DD] =  8'h20;
		ram[15'h18DE] =  8'h28;
		ram[15'h18DF] =  8'h3C;
		ram[15'h18E0] =  8'h69;
		ram[15'h18E1] =  8'h78;
		ram[15'h18E2] =  8'h2C;
		ram[15'h18E3] =  8'h69;
		ram[15'h18E4] =  8'h79;
		ram[15'h18E5] =  8'h3E;
		ram[15'h18E6] =  8'h2B;
		ram[15'h18E7] =  8'h31;
		ram[15'h18E8] =  8'h29;
		ram[15'h18E9] =  8'h2C;
		ram[15'h18EA] =  8'h3C;
		ram[15'h18EB] =  8'h62;
		ram[15'h18EC] =  8'h2C;
		ram[15'h18ED] =  8'h63;
		ram[15'h18EE] =  8'h2C;
		ram[15'h18EF] =  8'h64;
		ram[15'h18F0] =  8'h2C;
		ram[15'h18F1] =  8'h65;
		ram[15'h18F2] =  8'h3E;
		ram[15'h18F3] =  8'h2E;
		ram[15'h18F4] =  8'h2E;
		ram[15'h18F5] =  8'h2E;
		ram[15'h18F6] =  8'h2E;
		ram[15'h18F7] =  8'h2E;
		ram[15'h18F8] =  8'h2E;
		ram[15'h18F9] =  8'h24;
		ram[15'h18FA] =  8'hD7;
		ram[15'h18FB] =  8'hDD;
		ram[15'h18FC] =  8'h74;
		ram[15'h18FD] =  8'h01;
		ram[15'h18FE] =  8'h00;
		ram[15'h18FF] =  8'h64;
		ram[15'h1900] =  8'hB6;
		ram[15'h1901] =  8'h39;
		ram[15'h1902] =  8'h00;
		ram[15'h1903] =  8'h39;
		ram[15'h1904] =  8'h00;
		ram[15'h1905] =  8'hAC;
		ram[15'h1906] =  8'hE8;
		ram[15'h1907] =  8'hF5;
		ram[15'h1908] =  8'hB5;
		ram[15'h1909] =  8'hFE;
		ram[15'h190A] =  8'hAA;
		ram[15'h190B] =  8'h12;
		ram[15'h190C] =  8'h10;
		ram[15'h190D] =  8'h66;
		ram[15'h190E] =  8'h95;
		ram[15'h190F] =  8'h20;
		ram[15'h1910] =  8'h01;
		ram[15'h1911] =  8'h00;
		ram[15'h1912] =  8'h00;
		ram[15'h1913] =  8'h00;
		ram[15'h1914] =  8'h00;
		ram[15'h1915] =  8'h01;
		ram[15'h1916] =  8'h00;
		ram[15'h1917] =  8'h01;
		ram[15'h1918] =  8'h00;
		ram[15'h1919] =  8'h00;
		ram[15'h191A] =  8'h00;
		ram[15'h191B] =  8'h00;
		ram[15'h191C] =  8'h00;
		ram[15'h191D] =  8'h00;
		ram[15'h191E] =  8'h00;
		ram[15'h191F] =  8'h00;
		ram[15'h1920] =  8'h00;
		ram[15'h1921] =  8'h00;
		ram[15'h1922] =  8'h00;
		ram[15'h1923] =  8'h00;
		ram[15'h1924] =  8'h00;
		ram[15'h1925] =  8'h00;
		ram[15'h1926] =  8'h00;
		ram[15'h1927] =  8'h00;
		ram[15'h1928] =  8'h00;
		ram[15'h1929] =  8'h00;
		ram[15'h192A] =  8'h00;
		ram[15'h192B] =  8'h00;
		ram[15'h192C] =  8'h00;
		ram[15'h192D] =  8'hFF;
		ram[15'h192E] =  8'hFF;
		ram[15'h192F] =  8'h00;
		ram[15'h1930] =  8'h00;
		ram[15'h1931] =  8'h00;
		ram[15'h1932] =  8'h00;
		ram[15'h1933] =  8'h00;
		ram[15'h1934] =  8'h00;
		ram[15'h1935] =  8'h00;
		ram[15'h1936] =  8'h00;
		ram[15'h1937] =  8'h6A;
		ram[15'h1938] =  8'h1A;
		ram[15'h1939] =  8'h88;
		ram[15'h193A] =  8'h31;
		ram[15'h193B] =  8'h6C;
		ram[15'h193C] =  8'h64;
		ram[15'h193D] =  8'h20;
		ram[15'h193E] =  8'h28;
		ram[15'h193F] =  8'h3C;
		ram[15'h1940] =  8'h69;
		ram[15'h1941] =  8'h78;
		ram[15'h1942] =  8'h2C;
		ram[15'h1943] =  8'h69;
		ram[15'h1944] =  8'h79;
		ram[15'h1945] =  8'h3E;
		ram[15'h1946] =  8'h2B;
		ram[15'h1947] =  8'h31;
		ram[15'h1948] =  8'h29;
		ram[15'h1949] =  8'h2C;
		ram[15'h194A] =  8'h3C;
		ram[15'h194B] =  8'h68;
		ram[15'h194C] =  8'h2C;
		ram[15'h194D] =  8'h6C;
		ram[15'h194E] =  8'h3E;
		ram[15'h194F] =  8'h2E;
		ram[15'h1950] =  8'h2E;
		ram[15'h1951] =  8'h2E;
		ram[15'h1952] =  8'h2E;
		ram[15'h1953] =  8'h2E;
		ram[15'h1954] =  8'h2E;
		ram[15'h1955] =  8'h2E;
		ram[15'h1956] =  8'h2E;
		ram[15'h1957] =  8'h2E;
		ram[15'h1958] =  8'h2E;
		ram[15'h1959] =  8'h24;
		ram[15'h195A] =  8'hD7;
		ram[15'h195B] =  8'hDD;
		ram[15'h195C] =  8'h77;
		ram[15'h195D] =  8'h01;
		ram[15'h195E] =  8'h00;
		ram[15'h195F] =  8'hAF;
		ram[15'h1960] =  8'h67;
		ram[15'h1961] =  8'h39;
		ram[15'h1962] =  8'h00;
		ram[15'h1963] =  8'h39;
		ram[15'h1964] =  8'h00;
		ram[15'h1965] =  8'h13;
		ram[15'h1966] =  8'h4F;
		ram[15'h1967] =  8'h44;
		ram[15'h1968] =  8'h06;
		ram[15'h1969] =  8'hD7;
		ram[15'h196A] =  8'hBC;
		ram[15'h196B] =  8'h50;
		ram[15'h196C] =  8'hAC;
		ram[15'h196D] =  8'hAF;
		ram[15'h196E] =  8'h5F;
		ram[15'h196F] =  8'h20;
		ram[15'h1970] =  8'h00;
		ram[15'h1971] =  8'h00;
		ram[15'h1972] =  8'h00;
		ram[15'h1973] =  8'h00;
		ram[15'h1974] =  8'h00;
		ram[15'h1975] =  8'h01;
		ram[15'h1976] =  8'h00;
		ram[15'h1977] =  8'h01;
		ram[15'h1978] =  8'h00;
		ram[15'h1979] =  8'h00;
		ram[15'h197A] =  8'h00;
		ram[15'h197B] =  8'h00;
		ram[15'h197C] =  8'h00;
		ram[15'h197D] =  8'h00;
		ram[15'h197E] =  8'h00;
		ram[15'h197F] =  8'h00;
		ram[15'h1980] =  8'h00;
		ram[15'h1981] =  8'h00;
		ram[15'h1982] =  8'h00;
		ram[15'h1983] =  8'h00;
		ram[15'h1984] =  8'h00;
		ram[15'h1985] =  8'h00;
		ram[15'h1986] =  8'h00;
		ram[15'h1987] =  8'h00;
		ram[15'h1988] =  8'h00;
		ram[15'h1989] =  8'h00;
		ram[15'h198A] =  8'h00;
		ram[15'h198B] =  8'h00;
		ram[15'h198C] =  8'h00;
		ram[15'h198D] =  8'h00;
		ram[15'h198E] =  8'h00;
		ram[15'h198F] =  8'h00;
		ram[15'h1990] =  8'h00;
		ram[15'h1991] =  8'h00;
		ram[15'h1992] =  8'h00;
		ram[15'h1993] =  8'h00;
		ram[15'h1994] =  8'hFF;
		ram[15'h1995] =  8'h00;
		ram[15'h1996] =  8'h00;
		ram[15'h1997] =  8'hCC;
		ram[15'h1998] =  8'hBE;
		ram[15'h1999] =  8'h5A;
		ram[15'h199A] =  8'h96;
		ram[15'h199B] =  8'h6C;
		ram[15'h199C] =  8'h64;
		ram[15'h199D] =  8'h20;
		ram[15'h199E] =  8'h28;
		ram[15'h199F] =  8'h3C;
		ram[15'h19A0] =  8'h69;
		ram[15'h19A1] =  8'h78;
		ram[15'h19A2] =  8'h2C;
		ram[15'h19A3] =  8'h69;
		ram[15'h19A4] =  8'h79;
		ram[15'h19A5] =  8'h3E;
		ram[15'h19A6] =  8'h2B;
		ram[15'h19A7] =  8'h31;
		ram[15'h19A8] =  8'h29;
		ram[15'h19A9] =  8'h2C;
		ram[15'h19AA] =  8'h61;
		ram[15'h19AB] =  8'h2E;
		ram[15'h19AC] =  8'h2E;
		ram[15'h19AD] =  8'h2E;
		ram[15'h19AE] =  8'h2E;
		ram[15'h19AF] =  8'h2E;
		ram[15'h19B0] =  8'h2E;
		ram[15'h19B1] =  8'h2E;
		ram[15'h19B2] =  8'h2E;
		ram[15'h19B3] =  8'h2E;
		ram[15'h19B4] =  8'h2E;
		ram[15'h19B5] =  8'h2E;
		ram[15'h19B6] =  8'h2E;
		ram[15'h19B7] =  8'h2E;
		ram[15'h19B8] =  8'h2E;
		ram[15'h19B9] =  8'h24;
		ram[15'h19BA] =  8'hD7;
		ram[15'h19BB] =  8'h02;
		ram[15'h19BC] =  8'h00;
		ram[15'h19BD] =  8'h00;
		ram[15'h19BE] =  8'h00;
		ram[15'h19BF] =  8'h3B;
		ram[15'h19C0] =  8'h0C;
		ram[15'h19C1] =  8'h92;
		ram[15'h19C2] =  8'hB5;
		ram[15'h19C3] =  8'hFF;
		ram[15'h19C4] =  8'h6C;
		ram[15'h19C5] =  8'h9E;
		ram[15'h19C6] =  8'h95;
		ram[15'h19C7] =  8'h3A;
		ram[15'h19C8] =  8'h00;
		ram[15'h19C9] =  8'h3B;
		ram[15'h19CA] =  8'h00;
		ram[15'h19CB] =  8'hC1;
		ram[15'h19CC] =  8'h21;
		ram[15'h19CD] =  8'hE7;
		ram[15'h19CE] =  8'hBD;
		ram[15'h19CF] =  8'h18;
		ram[15'h19D0] =  8'h00;
		ram[15'h19D1] =  8'h00;
		ram[15'h19D2] =  8'h00;
		ram[15'h19D3] =  8'h00;
		ram[15'h19D4] =  8'h00;
		ram[15'h19D5] =  8'h00;
		ram[15'h19D6] =  8'h00;
		ram[15'h19D7] =  8'h00;
		ram[15'h19D8] =  8'h00;
		ram[15'h19D9] =  8'h00;
		ram[15'h19DA] =  8'h00;
		ram[15'h19DB] =  8'h00;
		ram[15'h19DC] =  8'h00;
		ram[15'h19DD] =  8'h00;
		ram[15'h19DE] =  8'h00;
		ram[15'h19DF] =  8'h00;
		ram[15'h19E0] =  8'h00;
		ram[15'h19E1] =  8'h00;
		ram[15'h19E2] =  8'h00;
		ram[15'h19E3] =  8'h00;
		ram[15'h19E4] =  8'h00;
		ram[15'h19E5] =  8'h00;
		ram[15'h19E6] =  8'h00;
		ram[15'h19E7] =  8'hFF;
		ram[15'h19E8] =  8'hFF;
		ram[15'h19E9] =  8'h00;
		ram[15'h19EA] =  8'h00;
		ram[15'h19EB] =  8'h00;
		ram[15'h19EC] =  8'h00;
		ram[15'h19ED] =  8'h00;
		ram[15'h19EE] =  8'h00;
		ram[15'h19EF] =  8'h00;
		ram[15'h19F0] =  8'h00;
		ram[15'h19F1] =  8'h00;
		ram[15'h19F2] =  8'h00;
		ram[15'h19F3] =  8'h00;
		ram[15'h19F4] =  8'hFF;
		ram[15'h19F5] =  8'h00;
		ram[15'h19F6] =  8'h00;
		ram[15'h19F7] =  8'h7A;
		ram[15'h19F8] =  8'h4C;
		ram[15'h19F9] =  8'h11;
		ram[15'h19FA] =  8'h4F;
		ram[15'h19FB] =  8'h6C;
		ram[15'h19FC] =  8'h64;
		ram[15'h19FD] =  8'h20;
		ram[15'h19FE] =  8'h28;
		ram[15'h19FF] =  8'h3C;
		ram[15'h1A00] =  8'h62;
		ram[15'h1A01] =  8'h63;
		ram[15'h1A02] =  8'h2C;
		ram[15'h1A03] =  8'h64;
		ram[15'h1A04] =  8'h65;
		ram[15'h1A05] =  8'h3E;
		ram[15'h1A06] =  8'h29;
		ram[15'h1A07] =  8'h2C;
		ram[15'h1A08] =  8'h61;
		ram[15'h1A09] =  8'h2E;
		ram[15'h1A0A] =  8'h2E;
		ram[15'h1A0B] =  8'h2E;
		ram[15'h1A0C] =  8'h2E;
		ram[15'h1A0D] =  8'h2E;
		ram[15'h1A0E] =  8'h2E;
		ram[15'h1A0F] =  8'h2E;
		ram[15'h1A10] =  8'h2E;
		ram[15'h1A11] =  8'h2E;
		ram[15'h1A12] =  8'h2E;
		ram[15'h1A13] =  8'h2E;
		ram[15'h1A14] =  8'h2E;
		ram[15'h1A15] =  8'h2E;
		ram[15'h1A16] =  8'h2E;
		ram[15'h1A17] =  8'h2E;
		ram[15'h1A18] =  8'h2E;
		ram[15'h1A19] =  8'h24;
		ram[15'h1A1A] =  8'hE5;
		ram[15'h1A1B] =  8'h7E;
		ram[15'h1A1C] =  8'h23;
		ram[15'h1A1D] =  8'h66;
		ram[15'h1A1E] =  8'h6F;
		ram[15'h1A1F] =  8'h7E;
		ram[15'h1A20] =  8'h32;
		ram[15'h1A21] =  8'hA3;
		ram[15'h1A22] =  8'h1C;
		ram[15'h1A23] =  8'h23;
		ram[15'h1A24] =  8'hE5;
		ram[15'h1A25] =  8'h11;
		ram[15'h1A26] =  8'h14;
		ram[15'h1A27] =  8'h00;
		ram[15'h1A28] =  8'h19;
		ram[15'h1A29] =  8'h11;
		ram[15'h1A2A] =  8'h14;
		ram[15'h1A2B] =  8'h1C;
		ram[15'h1A2C] =  8'hCD;
		ram[15'h1A2D] =  8'h83;
		ram[15'h1A2E] =  8'h1B;
		ram[15'h1A2F] =  8'hE1;
		ram[15'h1A30] =  8'hE5;
		ram[15'h1A31] =  8'h11;
		ram[15'h1A32] =  8'h28;
		ram[15'h1A33] =  8'h00;
		ram[15'h1A34] =  8'h19;
		ram[15'h1A35] =  8'h11;
		ram[15'h1A36] =  8'h3C;
		ram[15'h1A37] =  8'h1C;
		ram[15'h1A38] =  8'hCD;
		ram[15'h1A39] =  8'h83;
		ram[15'h1A3A] =  8'h1B;
		ram[15'h1A3B] =  8'h21;
		ram[15'h1A3C] =  8'h3C;
		ram[15'h1A3D] =  8'h1C;
		ram[15'h1A3E] =  8'h36;
		ram[15'h1A3F] =  8'h01;
		ram[15'h1A40] =  8'hE1;
		ram[15'h1A41] =  8'hE5;
		ram[15'h1A42] =  8'h11;
		ram[15'h1A43] =  8'h7E;
		ram[15'h1A44] =  8'h1C;
		ram[15'h1A45] =  8'h01;
		ram[15'h1A46] =  8'h04;
		ram[15'h1A47] =  8'h00;
		ram[15'h1A48] =  8'hED;
		ram[15'h1A49] =  8'hB0;
		ram[15'h1A4A] =  8'h11;
		ram[15'h1A4B] =  8'h3A;
		ram[15'h1A4C] =  8'h00;
		ram[15'h1A4D] =  8'h01;
		ram[15'h1A4E] =  8'h10;
		ram[15'h1A4F] =  8'h00;
		ram[15'h1A50] =  8'hED;
		ram[15'h1A51] =  8'hB0;
		ram[15'h1A52] =  8'h11;
		ram[15'h1A53] =  8'h2C;
		ram[15'h1A54] =  8'h00;
		ram[15'h1A55] =  8'h19;
		ram[15'h1A56] =  8'hEB;
		ram[15'h1A57] =  8'h0E;
		ram[15'h1A58] =  8'h09;
		ram[15'h1A59] =  8'hCD;
		ram[15'h1A5A] =  8'h0C;
		ram[15'h1A5B] =  8'h1D;
		ram[15'h1A5C] =  8'hCD;
		ram[15'h1A5D] =  8'hBE;
		ram[15'h1A5E] =  8'h1D;
		ram[15'h1A5F] =  8'h3A;
		ram[15'h1A60] =  8'h7E;
		ram[15'h1A61] =  8'h1C;
		ram[15'h1A62] =  8'hFE;
		ram[15'h1A63] =  8'h76;
		ram[15'h1A64] =  8'hCA;
		ram[15'h1A65] =  8'h76;
		ram[15'h1A66] =  8'h1A;
		ram[15'h1A67] =  8'hE6;
		ram[15'h1A68] =  8'hDF;
		ram[15'h1A69] =  8'hFE;
		ram[15'h1A6A] =  8'hDD;
		ram[15'h1A6B] =  8'hC2;
		ram[15'h1A6C] =  8'h73;
		ram[15'h1A6D] =  8'h1A;
		ram[15'h1A6E] =  8'h3A;
		ram[15'h1A6F] =  8'h7F;
		ram[15'h1A70] =  8'h1C;
		ram[15'h1A71] =  8'hFE;
		ram[15'h1A72] =  8'h76;
		ram[15'h1A73] =  8'hC4;
		ram[15'h1A74] =  8'h64;
		ram[15'h1A75] =  8'h1C;
		ram[15'h1A76] =  8'hCD;
		ram[15'h1A77] =  8'hC3;
		ram[15'h1A78] =  8'h1B;
		ram[15'h1A79] =  8'hC4;
		ram[15'h1A7A] =  8'hE7;
		ram[15'h1A7B] =  8'h1B;
		ram[15'h1A7C] =  8'hE1;
		ram[15'h1A7D] =  8'hCA;
		ram[15'h1A7E] =  8'hB4;
		ram[15'h1A7F] =  8'h1A;
		ram[15'h1A80] =  8'h11;
		ram[15'h1A81] =  8'h3C;
		ram[15'h1A82] =  8'h00;
		ram[15'h1A83] =  8'h19;
		ram[15'h1A84] =  8'hCD;
		ram[15'h1A85] =  8'h7F;
		ram[15'h1A86] =  8'h1D;
		ram[15'h1A87] =  8'h11;
		ram[15'h1A88] =  8'h64;
		ram[15'h1A89] =  8'h1D;
		ram[15'h1A8A] =  8'hCA;
		ram[15'h1A8B] =  8'hAB;
		ram[15'h1A8C] =  8'h1A;
		ram[15'h1A8D] =  8'hE5;
		ram[15'h1A8E] =  8'h21;
		ram[15'h1A8F] =  8'hD2;
		ram[15'h1A90] =  8'h1D;
		ram[15'h1A91] =  8'h11;
		ram[15'h1A92] =  8'h69;
		ram[15'h1A93] =  8'h1D;
		ram[15'h1A94] =  8'h0E;
		ram[15'h1A95] =  8'h09;
		ram[15'h1A96] =  8'hCD;
		ram[15'h1A97] =  8'h0C;
		ram[15'h1A98] =  8'h1D;
		ram[15'h1A99] =  8'hCD;
		ram[15'h1A9A] =  8'hD7;
		ram[15'h1A9B] =  8'h1C;
		ram[15'h1A9C] =  8'h11;
		ram[15'h1A9D] =  8'h71;
		ram[15'h1A9E] =  8'h1D;
		ram[15'h1A9F] =  8'h0E;
		ram[15'h1AA0] =  8'h09;
		ram[15'h1AA1] =  8'hCD;
		ram[15'h1AA2] =  8'h0C;
		ram[15'h1AA3] =  8'h1D;
		ram[15'h1AA4] =  8'hE1;
		ram[15'h1AA5] =  8'hCD;
		ram[15'h1AA6] =  8'hD7;
		ram[15'h1AA7] =  8'h1C;
		ram[15'h1AA8] =  8'h11;
		ram[15'h1AA9] =  8'h7C;
		ram[15'h1AAA] =  8'h1D;
		ram[15'h1AAB] =  8'h0E;
		ram[15'h1AAC] =  8'h09;
		ram[15'h1AAD] =  8'hCD;
		ram[15'h1AAE] =  8'h0C;
		ram[15'h1AAF] =  8'h1D;
		ram[15'h1AB0] =  8'hE1;
		ram[15'h1AB1] =  8'h23;
		ram[15'h1AB2] =  8'h23;
		ram[15'h1AB3] =  8'hC9;
		ram[15'h1AB4] =  8'hE5;
		ram[15'h1AB5] =  8'h3E;
		ram[15'h1AB6] =  8'h01;
		ram[15'h1AB7] =  8'h32;
		ram[15'h1AB8] =  8'h2A;
		ram[15'h1AB9] =  8'h1B;
		ram[15'h1ABA] =  8'h32;
		ram[15'h1ABB] =  8'h4E;
		ram[15'h1ABC] =  8'h1B;
		ram[15'h1ABD] =  8'h21;
		ram[15'h1ABE] =  8'h14;
		ram[15'h1ABF] =  8'h1C;
		ram[15'h1AC0] =  8'h22;
		ram[15'h1AC1] =  8'h2B;
		ram[15'h1AC2] =  8'h1B;
		ram[15'h1AC3] =  8'h21;
		ram[15'h1AC4] =  8'h3C;
		ram[15'h1AC5] =  8'h1C;
		ram[15'h1AC6] =  8'h22;
		ram[15'h1AC7] =  8'h4F;
		ram[15'h1AC8] =  8'h1B;
		ram[15'h1AC9] =  8'h06;
		ram[15'h1ACA] =  8'h04;
		ram[15'h1ACB] =  8'hE1;
		ram[15'h1ACC] =  8'hE5;
		ram[15'h1ACD] =  8'h11;
		ram[15'h1ACE] =  8'h7E;
		ram[15'h1ACF] =  8'h1C;
		ram[15'h1AD0] =  8'hCD;
		ram[15'h1AD1] =  8'hDE;
		ram[15'h1AD2] =  8'h1A;
		ram[15'h1AD3] =  8'h06;
		ram[15'h1AD4] =  8'h10;
		ram[15'h1AD5] =  8'h11;
		ram[15'h1AD6] =  8'h3A;
		ram[15'h1AD7] =  8'h00;
		ram[15'h1AD8] =  8'hCD;
		ram[15'h1AD9] =  8'hDE;
		ram[15'h1ADA] =  8'h1A;
		ram[15'h1ADB] =  8'hC3;
		ram[15'h1ADC] =  8'h5F;
		ram[15'h1ADD] =  8'h1A;
		ram[15'h1ADE] =  8'hCD;
		ram[15'h1ADF] =  8'hE7;
		ram[15'h1AE0] =  8'h1A;
		ram[15'h1AE1] =  8'h23;
		ram[15'h1AE2] =  8'h05;
		ram[15'h1AE3] =  8'hC2;
		ram[15'h1AE4] =  8'hDE;
		ram[15'h1AE5] =  8'h1A;
		ram[15'h1AE6] =  8'hC9;
		ram[15'h1AE7] =  8'hC5;
		ram[15'h1AE8] =  8'hD5;
		ram[15'h1AE9] =  8'hE5;
		ram[15'h1AEA] =  8'h4E;
		ram[15'h1AEB] =  8'h11;
		ram[15'h1AEC] =  8'h14;
		ram[15'h1AED] =  8'h00;
		ram[15'h1AEE] =  8'h19;
		ram[15'h1AEF] =  8'h7E;
		ram[15'h1AF0] =  8'hFE;
		ram[15'h1AF1] =  8'h00;
		ram[15'h1AF2] =  8'hCA;
		ram[15'h1AF3] =  8'h08;
		ram[15'h1AF4] =  8'h1B;
		ram[15'h1AF5] =  8'h06;
		ram[15'h1AF6] =  8'h08;
		ram[15'h1AF7] =  8'h0F;
		ram[15'h1AF8] =  8'hF5;
		ram[15'h1AF9] =  8'h3E;
		ram[15'h1AFA] =  8'h00;
		ram[15'h1AFB] =  8'hDC;
		ram[15'h1AFC] =  8'h2D;
		ram[15'h1AFD] =  8'h1B;
		ram[15'h1AFE] =  8'hA9;
		ram[15'h1AFF] =  8'h0F;
		ram[15'h1B00] =  8'h4F;
		ram[15'h1B01] =  8'hF1;
		ram[15'h1B02] =  8'h05;
		ram[15'h1B03] =  8'hC2;
		ram[15'h1B04] =  8'hF7;
		ram[15'h1B05] =  8'h1A;
		ram[15'h1B06] =  8'h06;
		ram[15'h1B07] =  8'h08;
		ram[15'h1B08] =  8'h11;
		ram[15'h1B09] =  8'h14;
		ram[15'h1B0A] =  8'h00;
		ram[15'h1B0B] =  8'h19;
		ram[15'h1B0C] =  8'h7E;
		ram[15'h1B0D] =  8'hFE;
		ram[15'h1B0E] =  8'h00;
		ram[15'h1B0F] =  8'hCA;
		ram[15'h1B10] =  8'h23;
		ram[15'h1B11] =  8'h1B;
		ram[15'h1B12] =  8'h06;
		ram[15'h1B13] =  8'h08;
		ram[15'h1B14] =  8'h0F;
		ram[15'h1B15] =  8'hF5;
		ram[15'h1B16] =  8'h3E;
		ram[15'h1B17] =  8'h00;
		ram[15'h1B18] =  8'hDC;
		ram[15'h1B19] =  8'h51;
		ram[15'h1B1A] =  8'h1B;
		ram[15'h1B1B] =  8'hA9;
		ram[15'h1B1C] =  8'h0F;
		ram[15'h1B1D] =  8'h4F;
		ram[15'h1B1E] =  8'hF1;
		ram[15'h1B1F] =  8'h05;
		ram[15'h1B20] =  8'hC2;
		ram[15'h1B21] =  8'h14;
		ram[15'h1B22] =  8'h1B;
		ram[15'h1B23] =  8'hE1;
		ram[15'h1B24] =  8'hD1;
		ram[15'h1B25] =  8'h79;
		ram[15'h1B26] =  8'h12;
		ram[15'h1B27] =  8'h13;
		ram[15'h1B28] =  8'hC1;
		ram[15'h1B29] =  8'hC9;
		ram[15'h1B2A] =  8'h00;
		ram[15'h1B2B] =  8'h00;
		ram[15'h1B2C] =  8'h00;
		ram[15'h1B2D] =  8'hC5;
		ram[15'h1B2E] =  8'hE5;
		ram[15'h1B2F] =  8'h2A;
		ram[15'h1B30] =  8'h2B;
		ram[15'h1B31] =  8'h1B;
		ram[15'h1B32] =  8'h46;
		ram[15'h1B33] =  8'h21;
		ram[15'h1B34] =  8'h2A;
		ram[15'h1B35] =  8'h1B;
		ram[15'h1B36] =  8'h7E;
		ram[15'h1B37] =  8'h4F;
		ram[15'h1B38] =  8'h07;
		ram[15'h1B39] =  8'h77;
		ram[15'h1B3A] =  8'hFE;
		ram[15'h1B3B] =  8'h01;
		ram[15'h1B3C] =  8'hC2;
		ram[15'h1B3D] =  8'h46;
		ram[15'h1B3E] =  8'h1B;
		ram[15'h1B3F] =  8'h2A;
		ram[15'h1B40] =  8'h2B;
		ram[15'h1B41] =  8'h1B;
		ram[15'h1B42] =  8'h23;
		ram[15'h1B43] =  8'h22;
		ram[15'h1B44] =  8'h2B;
		ram[15'h1B45] =  8'h1B;
		ram[15'h1B46] =  8'h78;
		ram[15'h1B47] =  8'hA1;
		ram[15'h1B48] =  8'hE1;
		ram[15'h1B49] =  8'hC1;
		ram[15'h1B4A] =  8'hC8;
		ram[15'h1B4B] =  8'h3E;
		ram[15'h1B4C] =  8'h01;
		ram[15'h1B4D] =  8'hC9;
		ram[15'h1B4E] =  8'h00;
		ram[15'h1B4F] =  8'h00;
		ram[15'h1B50] =  8'h00;
		ram[15'h1B51] =  8'hC5;
		ram[15'h1B52] =  8'hE5;
		ram[15'h1B53] =  8'h2A;
		ram[15'h1B54] =  8'h4F;
		ram[15'h1B55] =  8'h1B;
		ram[15'h1B56] =  8'h46;
		ram[15'h1B57] =  8'h21;
		ram[15'h1B58] =  8'h4E;
		ram[15'h1B59] =  8'h1B;
		ram[15'h1B5A] =  8'h7E;
		ram[15'h1B5B] =  8'h4F;
		ram[15'h1B5C] =  8'h07;
		ram[15'h1B5D] =  8'h77;
		ram[15'h1B5E] =  8'hFE;
		ram[15'h1B5F] =  8'h01;
		ram[15'h1B60] =  8'hC2;
		ram[15'h1B61] =  8'h6A;
		ram[15'h1B62] =  8'h1B;
		ram[15'h1B63] =  8'h2A;
		ram[15'h1B64] =  8'h4F;
		ram[15'h1B65] =  8'h1B;
		ram[15'h1B66] =  8'h23;
		ram[15'h1B67] =  8'h22;
		ram[15'h1B68] =  8'h4F;
		ram[15'h1B69] =  8'h1B;
		ram[15'h1B6A] =  8'h78;
		ram[15'h1B6B] =  8'hA1;
		ram[15'h1B6C] =  8'hE1;
		ram[15'h1B6D] =  8'hC1;
		ram[15'h1B6E] =  8'hC8;
		ram[15'h1B6F] =  8'h3E;
		ram[15'h1B70] =  8'h01;
		ram[15'h1B71] =  8'hC9;
		ram[15'h1B72] =  8'hF5;
		ram[15'h1B73] =  8'hC5;
		ram[15'h1B74] =  8'hD5;
		ram[15'h1B75] =  8'hE5;
		ram[15'h1B76] =  8'h36;
		ram[15'h1B77] =  8'h00;
		ram[15'h1B78] =  8'h54;
		ram[15'h1B79] =  8'h5D;
		ram[15'h1B7A] =  8'h13;
		ram[15'h1B7B] =  8'h0B;
		ram[15'h1B7C] =  8'hED;
		ram[15'h1B7D] =  8'hB0;
		ram[15'h1B7E] =  8'hE1;
		ram[15'h1B7F] =  8'hD1;
		ram[15'h1B80] =  8'hC1;
		ram[15'h1B81] =  8'hF1;
		ram[15'h1B82] =  8'hC9;
		ram[15'h1B83] =  8'hD5;
		ram[15'h1B84] =  8'hEB;
		ram[15'h1B85] =  8'h01;
		ram[15'h1B86] =  8'h28;
		ram[15'h1B87] =  8'h00;
		ram[15'h1B88] =  8'hCD;
		ram[15'h1B89] =  8'h72;
		ram[15'h1B8A] =  8'h1B;
		ram[15'h1B8B] =  8'hEB;
		ram[15'h1B8C] =  8'h06;
		ram[15'h1B8D] =  8'h14;
		ram[15'h1B8E] =  8'h0E;
		ram[15'h1B8F] =  8'h01;
		ram[15'h1B90] =  8'h16;
		ram[15'h1B91] =  8'h00;
		ram[15'h1B92] =  8'h5E;
		ram[15'h1B93] =  8'h7B;
		ram[15'h1B94] =  8'hA1;
		ram[15'h1B95] =  8'hCA;
		ram[15'h1B96] =  8'h99;
		ram[15'h1B97] =  8'h1B;
		ram[15'h1B98] =  8'h14;
		ram[15'h1B99] =  8'h79;
		ram[15'h1B9A] =  8'h07;
		ram[15'h1B9B] =  8'h4F;
		ram[15'h1B9C] =  8'hFE;
		ram[15'h1B9D] =  8'h01;
		ram[15'h1B9E] =  8'hC2;
		ram[15'h1B9F] =  8'h93;
		ram[15'h1BA0] =  8'h1B;
		ram[15'h1BA1] =  8'h23;
		ram[15'h1BA2] =  8'h05;
		ram[15'h1BA3] =  8'hC2;
		ram[15'h1BA4] =  8'h92;
		ram[15'h1BA5] =  8'h1B;
		ram[15'h1BA6] =  8'h7A;
		ram[15'h1BA7] =  8'hE6;
		ram[15'h1BA8] =  8'hF8;
		ram[15'h1BA9] =  8'h0F;
		ram[15'h1BAA] =  8'h0F;
		ram[15'h1BAB] =  8'h0F;
		ram[15'h1BAC] =  8'h6F;
		ram[15'h1BAD] =  8'h26;
		ram[15'h1BAE] =  8'h00;
		ram[15'h1BAF] =  8'h7A;
		ram[15'h1BB0] =  8'hE6;
		ram[15'h1BB1] =  8'h07;
		ram[15'h1BB2] =  8'h3C;
		ram[15'h1BB3] =  8'h47;
		ram[15'h1BB4] =  8'h3E;
		ram[15'h1BB5] =  8'h80;
		ram[15'h1BB6] =  8'h07;
		ram[15'h1BB7] =  8'h05;
		ram[15'h1BB8] =  8'hC2;
		ram[15'h1BB9] =  8'hB6;
		ram[15'h1BBA] =  8'h1B;
		ram[15'h1BBB] =  8'hD1;
		ram[15'h1BBC] =  8'h19;
		ram[15'h1BBD] =  8'h11;
		ram[15'h1BBE] =  8'h14;
		ram[15'h1BBF] =  8'h00;
		ram[15'h1BC0] =  8'h19;
		ram[15'h1BC1] =  8'h77;
		ram[15'h1BC2] =  8'hC9;
		ram[15'h1BC3] =  8'hC5;
		ram[15'h1BC4] =  8'hD5;
		ram[15'h1BC5] =  8'hE5;
		ram[15'h1BC6] =  8'h21;
		ram[15'h1BC7] =  8'h14;
		ram[15'h1BC8] =  8'h1C;
		ram[15'h1BC9] =  8'h11;
		ram[15'h1BCA] =  8'h14;
		ram[15'h1BCB] =  8'h00;
		ram[15'h1BCC] =  8'hEB;
		ram[15'h1BCD] =  8'h19;
		ram[15'h1BCE] =  8'hEB;
		ram[15'h1BCF] =  8'h34;
		ram[15'h1BD0] =  8'h7E;
		ram[15'h1BD1] =  8'hFE;
		ram[15'h1BD2] =  8'h00;
		ram[15'h1BD3] =  8'hCA;
		ram[15'h1BD4] =  8'hE2;
		ram[15'h1BD5] =  8'h1B;
		ram[15'h1BD6] =  8'h47;
		ram[15'h1BD7] =  8'h1A;
		ram[15'h1BD8] =  8'hA0;
		ram[15'h1BD9] =  8'hCA;
		ram[15'h1BDA] =  8'hDE;
		ram[15'h1BDB] =  8'h1B;
		ram[15'h1BDC] =  8'h36;
		ram[15'h1BDD] =  8'h00;
		ram[15'h1BDE] =  8'hC1;
		ram[15'h1BDF] =  8'hD1;
		ram[15'h1BE0] =  8'hE1;
		ram[15'h1BE1] =  8'hC9;
		ram[15'h1BE2] =  8'h23;
		ram[15'h1BE3] =  8'h13;
		ram[15'h1BE4] =  8'hC3;
		ram[15'h1BE5] =  8'hCF;
		ram[15'h1BE6] =  8'h1B;
		ram[15'h1BE7] =  8'hC5;
		ram[15'h1BE8] =  8'hD5;
		ram[15'h1BE9] =  8'hE5;
		ram[15'h1BEA] =  8'h21;
		ram[15'h1BEB] =  8'h3C;
		ram[15'h1BEC] =  8'h1C;
		ram[15'h1BED] =  8'h11;
		ram[15'h1BEE] =  8'h14;
		ram[15'h1BEF] =  8'h00;
		ram[15'h1BF0] =  8'hEB;
		ram[15'h1BF1] =  8'h19;
		ram[15'h1BF2] =  8'hEB;
		ram[15'h1BF3] =  8'h7E;
		ram[15'h1BF4] =  8'hB7;
		ram[15'h1BF5] =  8'hCA;
		ram[15'h1BF6] =  8'h0F;
		ram[15'h1BF7] =  8'h1C;
		ram[15'h1BF8] =  8'h47;
		ram[15'h1BF9] =  8'h1A;
		ram[15'h1BFA] =  8'hA0;
		ram[15'h1BFB] =  8'hC2;
		ram[15'h1BFC] =  8'h0B;
		ram[15'h1BFD] =  8'h1C;
		ram[15'h1BFE] =  8'h78;
		ram[15'h1BFF] =  8'h07;
		ram[15'h1C00] =  8'hFE;
		ram[15'h1C01] =  8'h01;
		ram[15'h1C02] =  8'hC2;
		ram[15'h1C03] =  8'h09;
		ram[15'h1C04] =  8'h1C;
		ram[15'h1C05] =  8'h36;
		ram[15'h1C06] =  8'h00;
		ram[15'h1C07] =  8'h23;
		ram[15'h1C08] =  8'h13;
		ram[15'h1C09] =  8'h77;
		ram[15'h1C0A] =  8'hAF;
		ram[15'h1C0B] =  8'hE1;
		ram[15'h1C0C] =  8'hD1;
		ram[15'h1C0D] =  8'hC1;
		ram[15'h1C0E] =  8'hC9;
		ram[15'h1C0F] =  8'h23;
		ram[15'h1C10] =  8'h13;
		ram[15'h1C11] =  8'hC3;
		ram[15'h1C12] =  8'hF3;
		ram[15'h1C13] =  8'h1B;
		ram[15'h1C14] =  8'h00;
		ram[15'h1C15] =  8'h00;
		ram[15'h1C16] =  8'h00;
		ram[15'h1C17] =  8'h00;
		ram[15'h1C18] =  8'h00;
		ram[15'h1C19] =  8'h00;
		ram[15'h1C1A] =  8'h00;
		ram[15'h1C1B] =  8'h00;
		ram[15'h1C1C] =  8'h00;
		ram[15'h1C1D] =  8'h00;
		ram[15'h1C1E] =  8'h00;
		ram[15'h1C1F] =  8'h00;
		ram[15'h1C20] =  8'h00;
		ram[15'h1C21] =  8'h00;
		ram[15'h1C22] =  8'h00;
		ram[15'h1C23] =  8'h00;
		ram[15'h1C24] =  8'h00;
		ram[15'h1C25] =  8'h00;
		ram[15'h1C26] =  8'h00;
		ram[15'h1C27] =  8'h00;
		ram[15'h1C28] =  8'h00;
		ram[15'h1C29] =  8'h00;
		ram[15'h1C2A] =  8'h00;
		ram[15'h1C2B] =  8'h00;
		ram[15'h1C2C] =  8'h00;
		ram[15'h1C2D] =  8'h00;
		ram[15'h1C2E] =  8'h00;
		ram[15'h1C2F] =  8'h00;
		ram[15'h1C30] =  8'h00;
		ram[15'h1C31] =  8'h00;
		ram[15'h1C32] =  8'h00;
		ram[15'h1C33] =  8'h00;
		ram[15'h1C34] =  8'h00;
		ram[15'h1C35] =  8'h00;
		ram[15'h1C36] =  8'h00;
		ram[15'h1C37] =  8'h00;
		ram[15'h1C38] =  8'h00;
		ram[15'h1C39] =  8'h00;
		ram[15'h1C3A] =  8'h00;
		ram[15'h1C3B] =  8'h00;
		ram[15'h1C3C] =  8'h00;
		ram[15'h1C3D] =  8'h00;
		ram[15'h1C3E] =  8'h00;
		ram[15'h1C3F] =  8'h00;
		ram[15'h1C40] =  8'h00;
		ram[15'h1C41] =  8'h00;
		ram[15'h1C42] =  8'h00;
		ram[15'h1C43] =  8'h00;
		ram[15'h1C44] =  8'h00;
		ram[15'h1C45] =  8'h00;
		ram[15'h1C46] =  8'h00;
		ram[15'h1C47] =  8'h00;
		ram[15'h1C48] =  8'h00;
		ram[15'h1C49] =  8'h00;
		ram[15'h1C4A] =  8'h00;
		ram[15'h1C4B] =  8'h00;
		ram[15'h1C4C] =  8'h00;
		ram[15'h1C4D] =  8'h00;
		ram[15'h1C4E] =  8'h00;
		ram[15'h1C4F] =  8'h00;
		ram[15'h1C50] =  8'h00;
		ram[15'h1C51] =  8'h00;
		ram[15'h1C52] =  8'h00;
		ram[15'h1C53] =  8'h00;
		ram[15'h1C54] =  8'h00;
		ram[15'h1C55] =  8'h00;
		ram[15'h1C56] =  8'h00;
		ram[15'h1C57] =  8'h00;
		ram[15'h1C58] =  8'h00;
		ram[15'h1C59] =  8'h00;
		ram[15'h1C5A] =  8'h00;
		ram[15'h1C5B] =  8'h00;
		ram[15'h1C5C] =  8'h00;
		ram[15'h1C5D] =  8'h00;
		ram[15'h1C5E] =  8'h00;
		ram[15'h1C5F] =  8'h00;
		ram[15'h1C60] =  8'h00;
		ram[15'h1C61] =  8'h00;
		ram[15'h1C62] =  8'h00;
		ram[15'h1C63] =  8'h00;
		ram[15'h1C64] =  8'hF5;
		ram[15'h1C65] =  8'hC5;
		ram[15'h1C66] =  8'hD5;
		ram[15'h1C67] =  8'hE5;
		ram[15'h1C68] =  8'hFD;
		ram[15'h1C69] =  8'hE5;
		ram[15'h1C6A] =  8'hF3;
		ram[15'h1C6B] =  8'hED;
		ram[15'h1C6C] =  8'h73;
		ram[15'h1C6D] =  8'hCB;
		ram[15'h1C6E] =  8'h1C;
		ram[15'h1C6F] =  8'h31;
		ram[15'h1C70] =  8'h3C;
		ram[15'h1C71] =  8'h00;
		ram[15'h1C72] =  8'hFD;
		ram[15'h1C73] =  8'hE1;
		ram[15'h1C74] =  8'hDD;
		ram[15'h1C75] =  8'hE1;
		ram[15'h1C76] =  8'hE1;
		ram[15'h1C77] =  8'hD1;
		ram[15'h1C78] =  8'hC1;
		ram[15'h1C79] =  8'hF1;
		ram[15'h1C7A] =  8'hED;
		ram[15'h1C7B] =  8'h7B;
		ram[15'h1C7C] =  8'h48;
		ram[15'h1C7D] =  8'h00;
		ram[15'h1C7E] =  8'h00;
		ram[15'h1C7F] =  8'h00;
		ram[15'h1C80] =  8'h00;
		ram[15'h1C81] =  8'h00;
		ram[15'h1C82] =  8'hED;
		ram[15'h1C83] =  8'h73;
		ram[15'h1C84] =  8'hC9;
		ram[15'h1C85] =  8'h1C;
		ram[15'h1C86] =  8'h31;
		ram[15'h1C87] =  8'hC9;
		ram[15'h1C88] =  8'h1C;
		ram[15'h1C89] =  8'hF5;
		ram[15'h1C8A] =  8'hC5;
		ram[15'h1C8B] =  8'hD5;
		ram[15'h1C8C] =  8'hE5;
		ram[15'h1C8D] =  8'hDD;
		ram[15'h1C8E] =  8'hE5;
		ram[15'h1C8F] =  8'hFD;
		ram[15'h1C90] =  8'hE5;
		ram[15'h1C91] =  8'hED;
		ram[15'h1C92] =  8'h7B;
		ram[15'h1C93] =  8'hCB;
		ram[15'h1C94] =  8'h1C;
		ram[15'h1C95] =  8'hFD;
		ram[15'h1C96] =  8'hE1;
		ram[15'h1C97] =  8'hFB;
		ram[15'h1C98] =  8'h2A;
		ram[15'h1C99] =  8'h3A;
		ram[15'h1C9A] =  8'h00;
		ram[15'h1C9B] =  8'h22;
		ram[15'h1C9C] =  8'hBB;
		ram[15'h1C9D] =  8'h1C;
		ram[15'h1C9E] =  8'h21;
		ram[15'h1C9F] =  8'hC7;
		ram[15'h1CA0] =  8'h1C;
		ram[15'h1CA1] =  8'h7E;
		ram[15'h1CA2] =  8'hE6;
		ram[15'h1CA3] =  8'hD7;
		ram[15'h1CA4] =  8'h77;
		ram[15'h1CA5] =  8'h06;
		ram[15'h1CA6] =  8'h10;
		ram[15'h1CA7] =  8'h11;
		ram[15'h1CA8] =  8'hBB;
		ram[15'h1CA9] =  8'h1C;
		ram[15'h1CAA] =  8'h21;
		ram[15'h1CAB] =  8'hD2;
		ram[15'h1CAC] =  8'h1D;
		ram[15'h1CAD] =  8'h1A;
		ram[15'h1CAE] =  8'h13;
		ram[15'h1CAF] =  8'hCD;
		ram[15'h1CB0] =  8'h96;
		ram[15'h1CB1] =  8'h1D;
		ram[15'h1CB2] =  8'h05;
		ram[15'h1CB3] =  8'hC2;
		ram[15'h1CB4] =  8'hAD;
		ram[15'h1CB5] =  8'h1C;
		ram[15'h1CB6] =  8'hE1;
		ram[15'h1CB7] =  8'hD1;
		ram[15'h1CB8] =  8'hC1;
		ram[15'h1CB9] =  8'hF1;
		ram[15'h1CBA] =  8'hC9;
		ram[15'h1CBB] =  8'h00;
		ram[15'h1CBC] =  8'h00;
		ram[15'h1CBD] =  8'h00;
		ram[15'h1CBE] =  8'h00;
		ram[15'h1CBF] =  8'h00;
		ram[15'h1CC0] =  8'h00;
		ram[15'h1CC1] =  8'h00;
		ram[15'h1CC2] =  8'h00;
		ram[15'h1CC3] =  8'h00;
		ram[15'h1CC4] =  8'h00;
		ram[15'h1CC5] =  8'h00;
		ram[15'h1CC6] =  8'h00;
		ram[15'h1CC7] =  8'h00;
		ram[15'h1CC8] =  8'h00;
		ram[15'h1CC9] =  8'h00;
		ram[15'h1CCA] =  8'h00;
		ram[15'h1CCB] =  8'h00;
		ram[15'h1CCC] =  8'h00;
		ram[15'h1CCD] =  8'h7E;
		ram[15'h1CCE] =  8'hCD;
		ram[15'h1CCF] =  8'hE9;
		ram[15'h1CD0] =  8'h1C;
		ram[15'h1CD1] =  8'h23;
		ram[15'h1CD2] =  8'h05;
		ram[15'h1CD3] =  8'hC2;
		ram[15'h1CD4] =  8'hCD;
		ram[15'h1CD5] =  8'h1C;
		ram[15'h1CD6] =  8'hC9;
		ram[15'h1CD7] =  8'hF5;
		ram[15'h1CD8] =  8'hC5;
		ram[15'h1CD9] =  8'hE5;
		ram[15'h1CDA] =  8'h06;
		ram[15'h1CDB] =  8'h04;
		ram[15'h1CDC] =  8'h7E;
		ram[15'h1CDD] =  8'hCD;
		ram[15'h1CDE] =  8'hE9;
		ram[15'h1CDF] =  8'h1C;
		ram[15'h1CE0] =  8'h23;
		ram[15'h1CE1] =  8'h05;
		ram[15'h1CE2] =  8'hC2;
		ram[15'h1CE3] =  8'hDC;
		ram[15'h1CE4] =  8'h1C;
		ram[15'h1CE5] =  8'hE1;
		ram[15'h1CE6] =  8'hC1;
		ram[15'h1CE7] =  8'hF1;
		ram[15'h1CE8] =  8'hC9;
		ram[15'h1CE9] =  8'hF5;
		ram[15'h1CEA] =  8'h0F;
		ram[15'h1CEB] =  8'h0F;
		ram[15'h1CEC] =  8'h0F;
		ram[15'h1CED] =  8'h0F;
		ram[15'h1CEE] =  8'hCD;
		ram[15'h1CEF] =  8'hF2;
		ram[15'h1CF0] =  8'h1C;
		ram[15'h1CF1] =  8'hF1;
		ram[15'h1CF2] =  8'hF5;
		ram[15'h1CF3] =  8'hC5;
		ram[15'h1CF4] =  8'hD5;
		ram[15'h1CF5] =  8'hE5;
		ram[15'h1CF6] =  8'hE6;
		ram[15'h1CF7] =  8'h0F;
		ram[15'h1CF8] =  8'hFE;
		ram[15'h1CF9] =  8'h0A;
		ram[15'h1CFA] =  8'hDA;
		ram[15'h1CFB] =  8'hFF;
		ram[15'h1CFC] =  8'h1C;
		ram[15'h1CFD] =  8'hC6;
		ram[15'h1CFE] =  8'h27;
		ram[15'h1CFF] =  8'hC6;
		ram[15'h1D00] =  8'h30;
		ram[15'h1D01] =  8'h5F;
		ram[15'h1D02] =  8'h0E;
		ram[15'h1D03] =  8'h02;
		ram[15'h1D04] =  8'hCD;
		ram[15'h1D05] =  8'h0C;
		ram[15'h1D06] =  8'h1D;
		ram[15'h1D07] =  8'hE1;
		ram[15'h1D08] =  8'hD1;
		ram[15'h1D09] =  8'hC1;
		ram[15'h1D0A] =  8'hF1;
		ram[15'h1D0B] =  8'hC9;
		ram[15'h1D0C] =  8'hF5;
		ram[15'h1D0D] =  8'hC5;
		ram[15'h1D0E] =  8'hD5;
		ram[15'h1D0F] =  8'hE5;
		ram[15'h1D10] =  8'h47;
		ram[15'h1D11] =  8'h79;
		ram[15'h1D12] =  8'hFE;
		ram[15'h1D13] =  8'h02;
		ram[15'h1D14] =  8'h28;
		ram[15'h1D15] =  8'h09;
		ram[15'h1D16] =  8'hFE;
		ram[15'h1D17] =  8'h09;
		ram[15'h1D18] =  8'h28;
		ram[15'h1D19] =  8'h0D;
		ram[15'h1D1A] =  8'hE1;
		ram[15'h1D1B] =  8'hD1;
		ram[15'h1D1C] =  8'hC1;
		ram[15'h1D1D] =  8'hF1;
		ram[15'h1D1E] =  8'hC9;
		ram[15'h1D1F] =  8'h78;
		ram[15'h1D20] =  8'hFE;
		ram[15'h1D21] =  8'h0A;
		ram[15'h1D22] =  8'h28;
		ram[15'h1D23] =  8'hF6;
		ram[15'h1D24] =  8'hD7;
		ram[15'h1D25] =  8'h18;
		ram[15'h1D26] =  8'hF3;
		ram[15'h1D27] =  8'h1A;
		ram[15'h1D28] =  8'hFE;
		ram[15'h1D29] =  8'h24;
		ram[15'h1D2A] =  8'h28;
		ram[15'h1D2B] =  8'hEE;
		ram[15'h1D2C] =  8'hFE;
		ram[15'h1D2D] =  8'h0A;
		ram[15'h1D2E] =  8'hC4;
		ram[15'h1D2F] =  8'h10;
		ram[15'h1D30] =  8'h00;
		ram[15'h1D31] =  8'h13;
		ram[15'h1D32] =  8'h18;
		ram[15'h1D33] =  8'hF3;
		ram[15'h1D34] =  8'h5A;
		ram[15'h1D35] =  8'h38;
		ram[15'h1D36] =  8'h30;
		ram[15'h1D37] =  8'h64;
		ram[15'h1D38] =  8'h6F;
		ram[15'h1D39] =  8'h63;
		ram[15'h1D3A] =  8'h20;
		ram[15'h1D3B] =  8'h69;
		ram[15'h1D3C] =  8'h6E;
		ram[15'h1D3D] =  8'h73;
		ram[15'h1D3E] =  8'h74;
		ram[15'h1D3F] =  8'h72;
		ram[15'h1D40] =  8'h75;
		ram[15'h1D41] =  8'h63;
		ram[15'h1D42] =  8'h74;
		ram[15'h1D43] =  8'h69;
		ram[15'h1D44] =  8'h6F;
		ram[15'h1D45] =  8'h6E;
		ram[15'h1D46] =  8'h20;
		ram[15'h1D47] =  8'h65;
		ram[15'h1D48] =  8'h78;
		ram[15'h1D49] =  8'h65;
		ram[15'h1D4A] =  8'h72;
		ram[15'h1D4B] =  8'h63;
		ram[15'h1D4C] =  8'h69;
		ram[15'h1D4D] =  8'h73;
		ram[15'h1D4E] =  8'h65;
		ram[15'h1D4F] =  8'h72;
		ram[15'h1D50] =  8'h0A;
		ram[15'h1D51] =  8'h0D;
		ram[15'h1D52] =  8'h0A;
		ram[15'h1D53] =  8'h0D;
		ram[15'h1D54] =  8'h24;
		ram[15'h1D55] =  8'h54;
		ram[15'h1D56] =  8'h65;
		ram[15'h1D57] =  8'h73;
		ram[15'h1D58] =  8'h74;
		ram[15'h1D59] =  8'h73;
		ram[15'h1D5A] =  8'h20;
		ram[15'h1D5B] =  8'h63;
		ram[15'h1D5C] =  8'h6F;
		ram[15'h1D5D] =  8'h6D;
		ram[15'h1D5E] =  8'h70;
		ram[15'h1D5F] =  8'h6C;
		ram[15'h1D60] =  8'h65;
		ram[15'h1D61] =  8'h74;
		ram[15'h1D62] =  8'h65;
		ram[15'h1D63] =  8'h24;
		ram[15'h1D64] =  8'h4F;
		ram[15'h1D65] =  8'h4B;
		ram[15'h1D66] =  8'h0A;
		ram[15'h1D67] =  8'h0D;
		ram[15'h1D68] =  8'h24;
		ram[15'h1D69] =  8'h20;
		ram[15'h1D6A] =  8'h20;
		ram[15'h1D6B] =  8'h20;
		ram[15'h1D6C] =  8'h43;
		ram[15'h1D6D] =  8'h52;
		ram[15'h1D6E] =  8'h43;
		ram[15'h1D6F] =  8'h3A;
		ram[15'h1D70] =  8'h24;
		ram[15'h1D71] =  8'h20;
		ram[15'h1D72] =  8'h65;
		ram[15'h1D73] =  8'h78;
		ram[15'h1D74] =  8'h70;
		ram[15'h1D75] =  8'h65;
		ram[15'h1D76] =  8'h63;
		ram[15'h1D77] =  8'h74;
		ram[15'h1D78] =  8'h65;
		ram[15'h1D79] =  8'h64;
		ram[15'h1D7A] =  8'h3A;
		ram[15'h1D7B] =  8'h24;
		ram[15'h1D7C] =  8'h0A;
		ram[15'h1D7D] =  8'h0D;
		ram[15'h1D7E] =  8'h24;
		ram[15'h1D7F] =  8'hC5;
		ram[15'h1D80] =  8'hD5;
		ram[15'h1D81] =  8'hE5;
		ram[15'h1D82] =  8'h11;
		ram[15'h1D83] =  8'hD2;
		ram[15'h1D84] =  8'h1D;
		ram[15'h1D85] =  8'h06;
		ram[15'h1D86] =  8'h04;
		ram[15'h1D87] =  8'h1A;
		ram[15'h1D88] =  8'hBE;
		ram[15'h1D89] =  8'hC2;
		ram[15'h1D8A] =  8'h92;
		ram[15'h1D8B] =  8'h1D;
		ram[15'h1D8C] =  8'h23;
		ram[15'h1D8D] =  8'h13;
		ram[15'h1D8E] =  8'h05;
		ram[15'h1D8F] =  8'hC2;
		ram[15'h1D90] =  8'h87;
		ram[15'h1D91] =  8'h1D;
		ram[15'h1D92] =  8'hE1;
		ram[15'h1D93] =  8'hD1;
		ram[15'h1D94] =  8'hC1;
		ram[15'h1D95] =  8'hC9;
		ram[15'h1D96] =  8'hF5;
		ram[15'h1D97] =  8'hC5;
		ram[15'h1D98] =  8'hD5;
		ram[15'h1D99] =  8'hE5;
		ram[15'h1D9A] =  8'hE5;
		ram[15'h1D9B] =  8'h11;
		ram[15'h1D9C] =  8'h03;
		ram[15'h1D9D] =  8'h00;
		ram[15'h1D9E] =  8'h19;
		ram[15'h1D9F] =  8'hAE;
		ram[15'h1DA0] =  8'h6F;
		ram[15'h1DA1] =  8'h26;
		ram[15'h1DA2] =  8'h00;
		ram[15'h1DA3] =  8'h29;
		ram[15'h1DA4] =  8'h29;
		ram[15'h1DA5] =  8'hEB;
		ram[15'h1DA6] =  8'h21;
		ram[15'h1DA7] =  8'hD6;
		ram[15'h1DA8] =  8'h1D;
		ram[15'h1DA9] =  8'h19;
		ram[15'h1DAA] =  8'hEB;
		ram[15'h1DAB] =  8'hE1;
		ram[15'h1DAC] =  8'h01;
		ram[15'h1DAD] =  8'h04;
		ram[15'h1DAE] =  8'h00;
		ram[15'h1DAF] =  8'h1A;
		ram[15'h1DB0] =  8'hA8;
		ram[15'h1DB1] =  8'h46;
		ram[15'h1DB2] =  8'h77;
		ram[15'h1DB3] =  8'h13;
		ram[15'h1DB4] =  8'h23;
		ram[15'h1DB5] =  8'h0D;
		ram[15'h1DB6] =  8'hC2;
		ram[15'h1DB7] =  8'hAF;
		ram[15'h1DB8] =  8'h1D;
		ram[15'h1DB9] =  8'hE1;
		ram[15'h1DBA] =  8'hD1;
		ram[15'h1DBB] =  8'hC1;
		ram[15'h1DBC] =  8'hF1;
		ram[15'h1DBD] =  8'hC9;
		ram[15'h1DBE] =  8'hF5;
		ram[15'h1DBF] =  8'hC5;
		ram[15'h1DC0] =  8'hE5;
		ram[15'h1DC1] =  8'h21;
		ram[15'h1DC2] =  8'hD2;
		ram[15'h1DC3] =  8'h1D;
		ram[15'h1DC4] =  8'h3E;
		ram[15'h1DC5] =  8'hFF;
		ram[15'h1DC6] =  8'h06;
		ram[15'h1DC7] =  8'h04;
		ram[15'h1DC8] =  8'h77;
		ram[15'h1DC9] =  8'h23;
		ram[15'h1DCA] =  8'h05;
		ram[15'h1DCB] =  8'hC2;
		ram[15'h1DCC] =  8'hC8;
		ram[15'h1DCD] =  8'h1D;
		ram[15'h1DCE] =  8'hE1;
		ram[15'h1DCF] =  8'hC1;
		ram[15'h1DD0] =  8'hF1;
		ram[15'h1DD1] =  8'hC9;
		ram[15'h1DD2] =  8'h00;
		ram[15'h1DD3] =  8'h00;
		ram[15'h1DD4] =  8'h00;
		ram[15'h1DD5] =  8'h00;
		ram[15'h1DD6] =  8'h00;
		ram[15'h1DD7] =  8'h00;
		ram[15'h1DD8] =  8'h00;
		ram[15'h1DD9] =  8'h00;
		ram[15'h1DDA] =  8'h77;
		ram[15'h1DDB] =  8'h07;
		ram[15'h1DDC] =  8'h30;
		ram[15'h1DDD] =  8'h96;
		ram[15'h1DDE] =  8'hEE;
		ram[15'h1DDF] =  8'h0E;
		ram[15'h1DE0] =  8'h61;
		ram[15'h1DE1] =  8'h2C;
		ram[15'h1DE2] =  8'h99;
		ram[15'h1DE3] =  8'h09;
		ram[15'h1DE4] =  8'h51;
		ram[15'h1DE5] =  8'hBA;
		ram[15'h1DE6] =  8'h07;
		ram[15'h1DE7] =  8'h6D;
		ram[15'h1DE8] =  8'hC4;
		ram[15'h1DE9] =  8'h19;
		ram[15'h1DEA] =  8'h70;
		ram[15'h1DEB] =  8'h6A;
		ram[15'h1DEC] =  8'hF4;
		ram[15'h1DED] =  8'h8F;
		ram[15'h1DEE] =  8'hE9;
		ram[15'h1DEF] =  8'h63;
		ram[15'h1DF0] =  8'hA5;
		ram[15'h1DF1] =  8'h35;
		ram[15'h1DF2] =  8'h9E;
		ram[15'h1DF3] =  8'h64;
		ram[15'h1DF4] =  8'h95;
		ram[15'h1DF5] =  8'hA3;
		ram[15'h1DF6] =  8'h0E;
		ram[15'h1DF7] =  8'hDB;
		ram[15'h1DF8] =  8'h88;
		ram[15'h1DF9] =  8'h32;
		ram[15'h1DFA] =  8'h79;
		ram[15'h1DFB] =  8'hDC;
		ram[15'h1DFC] =  8'hB8;
		ram[15'h1DFD] =  8'hA4;
		ram[15'h1DFE] =  8'hE0;
		ram[15'h1DFF] =  8'hD5;
		ram[15'h1E00] =  8'hE9;
		ram[15'h1E01] =  8'h1E;
		ram[15'h1E02] =  8'h97;
		ram[15'h1E03] =  8'hD2;
		ram[15'h1E04] =  8'hD9;
		ram[15'h1E05] =  8'h88;
		ram[15'h1E06] =  8'h09;
		ram[15'h1E07] =  8'hB6;
		ram[15'h1E08] =  8'h4C;
		ram[15'h1E09] =  8'h2B;
		ram[15'h1E0A] =  8'h7E;
		ram[15'h1E0B] =  8'hB1;
		ram[15'h1E0C] =  8'h7C;
		ram[15'h1E0D] =  8'hBD;
		ram[15'h1E0E] =  8'hE7;
		ram[15'h1E0F] =  8'hB8;
		ram[15'h1E10] =  8'h2D;
		ram[15'h1E11] =  8'h07;
		ram[15'h1E12] =  8'h90;
		ram[15'h1E13] =  8'hBF;
		ram[15'h1E14] =  8'h1D;
		ram[15'h1E15] =  8'h91;
		ram[15'h1E16] =  8'h1D;
		ram[15'h1E17] =  8'hB7;
		ram[15'h1E18] =  8'h10;
		ram[15'h1E19] =  8'h64;
		ram[15'h1E1A] =  8'h6A;
		ram[15'h1E1B] =  8'hB0;
		ram[15'h1E1C] =  8'h20;
		ram[15'h1E1D] =  8'hF2;
		ram[15'h1E1E] =  8'hF3;
		ram[15'h1E1F] =  8'hB9;
		ram[15'h1E20] =  8'h71;
		ram[15'h1E21] =  8'h48;
		ram[15'h1E22] =  8'h84;
		ram[15'h1E23] =  8'hBE;
		ram[15'h1E24] =  8'h41;
		ram[15'h1E25] =  8'hDE;
		ram[15'h1E26] =  8'h1A;
		ram[15'h1E27] =  8'hDA;
		ram[15'h1E28] =  8'hD4;
		ram[15'h1E29] =  8'h7D;
		ram[15'h1E2A] =  8'h6D;
		ram[15'h1E2B] =  8'hDD;
		ram[15'h1E2C] =  8'hE4;
		ram[15'h1E2D] =  8'hEB;
		ram[15'h1E2E] =  8'hF4;
		ram[15'h1E2F] =  8'hD4;
		ram[15'h1E30] =  8'hB5;
		ram[15'h1E31] =  8'h51;
		ram[15'h1E32] =  8'h83;
		ram[15'h1E33] =  8'hD3;
		ram[15'h1E34] =  8'h85;
		ram[15'h1E35] =  8'hC7;
		ram[15'h1E36] =  8'h13;
		ram[15'h1E37] =  8'h6C;
		ram[15'h1E38] =  8'h98;
		ram[15'h1E39] =  8'h56;
		ram[15'h1E3A] =  8'h64;
		ram[15'h1E3B] =  8'h6B;
		ram[15'h1E3C] =  8'hA8;
		ram[15'h1E3D] =  8'hC0;
		ram[15'h1E3E] =  8'hFD;
		ram[15'h1E3F] =  8'h62;
		ram[15'h1E40] =  8'hF9;
		ram[15'h1E41] =  8'h7A;
		ram[15'h1E42] =  8'h8A;
		ram[15'h1E43] =  8'h65;
		ram[15'h1E44] =  8'hC9;
		ram[15'h1E45] =  8'hEC;
		ram[15'h1E46] =  8'h14;
		ram[15'h1E47] =  8'h01;
		ram[15'h1E48] =  8'h5C;
		ram[15'h1E49] =  8'h4F;
		ram[15'h1E4A] =  8'h63;
		ram[15'h1E4B] =  8'h06;
		ram[15'h1E4C] =  8'h6C;
		ram[15'h1E4D] =  8'hD9;
		ram[15'h1E4E] =  8'hFA;
		ram[15'h1E4F] =  8'h0F;
		ram[15'h1E50] =  8'h3D;
		ram[15'h1E51] =  8'h63;
		ram[15'h1E52] =  8'h8D;
		ram[15'h1E53] =  8'h08;
		ram[15'h1E54] =  8'h0D;
		ram[15'h1E55] =  8'hF5;
		ram[15'h1E56] =  8'h3B;
		ram[15'h1E57] =  8'h6E;
		ram[15'h1E58] =  8'h20;
		ram[15'h1E59] =  8'hC8;
		ram[15'h1E5A] =  8'h4C;
		ram[15'h1E5B] =  8'h69;
		ram[15'h1E5C] =  8'h10;
		ram[15'h1E5D] =  8'h5E;
		ram[15'h1E5E] =  8'hD5;
		ram[15'h1E5F] =  8'h60;
		ram[15'h1E60] =  8'h41;
		ram[15'h1E61] =  8'hE4;
		ram[15'h1E62] =  8'hA2;
		ram[15'h1E63] =  8'h67;
		ram[15'h1E64] =  8'h71;
		ram[15'h1E65] =  8'h72;
		ram[15'h1E66] =  8'h3C;
		ram[15'h1E67] =  8'h03;
		ram[15'h1E68] =  8'hE4;
		ram[15'h1E69] =  8'hD1;
		ram[15'h1E6A] =  8'h4B;
		ram[15'h1E6B] =  8'h04;
		ram[15'h1E6C] =  8'hD4;
		ram[15'h1E6D] =  8'h47;
		ram[15'h1E6E] =  8'hD2;
		ram[15'h1E6F] =  8'h0D;
		ram[15'h1E70] =  8'h85;
		ram[15'h1E71] =  8'hFD;
		ram[15'h1E72] =  8'hA5;
		ram[15'h1E73] =  8'h0A;
		ram[15'h1E74] =  8'hB5;
		ram[15'h1E75] =  8'h6B;
		ram[15'h1E76] =  8'h35;
		ram[15'h1E77] =  8'hB5;
		ram[15'h1E78] =  8'hA8;
		ram[15'h1E79] =  8'hFA;
		ram[15'h1E7A] =  8'h42;
		ram[15'h1E7B] =  8'hB2;
		ram[15'h1E7C] =  8'h98;
		ram[15'h1E7D] =  8'h6C;
		ram[15'h1E7E] =  8'hDB;
		ram[15'h1E7F] =  8'hBB;
		ram[15'h1E80] =  8'hC9;
		ram[15'h1E81] =  8'hD6;
		ram[15'h1E82] =  8'hAC;
		ram[15'h1E83] =  8'hBC;
		ram[15'h1E84] =  8'hF9;
		ram[15'h1E85] =  8'h40;
		ram[15'h1E86] =  8'h32;
		ram[15'h1E87] =  8'hD8;
		ram[15'h1E88] =  8'h6C;
		ram[15'h1E89] =  8'hE3;
		ram[15'h1E8A] =  8'h45;
		ram[15'h1E8B] =  8'hDF;
		ram[15'h1E8C] =  8'h5C;
		ram[15'h1E8D] =  8'h75;
		ram[15'h1E8E] =  8'hDC;
		ram[15'h1E8F] =  8'hD6;
		ram[15'h1E90] =  8'h0D;
		ram[15'h1E91] =  8'hCF;
		ram[15'h1E92] =  8'hAB;
		ram[15'h1E93] =  8'hD1;
		ram[15'h1E94] =  8'h3D;
		ram[15'h1E95] =  8'h59;
		ram[15'h1E96] =  8'h26;
		ram[15'h1E97] =  8'hD9;
		ram[15'h1E98] =  8'h30;
		ram[15'h1E99] =  8'hAC;
		ram[15'h1E9A] =  8'h51;
		ram[15'h1E9B] =  8'hDE;
		ram[15'h1E9C] =  8'h00;
		ram[15'h1E9D] =  8'h3A;
		ram[15'h1E9E] =  8'hC8;
		ram[15'h1E9F] =  8'hD7;
		ram[15'h1EA0] =  8'h51;
		ram[15'h1EA1] =  8'h80;
		ram[15'h1EA2] =  8'hBF;
		ram[15'h1EA3] =  8'hD0;
		ram[15'h1EA4] =  8'h61;
		ram[15'h1EA5] =  8'h16;
		ram[15'h1EA6] =  8'h21;
		ram[15'h1EA7] =  8'hB4;
		ram[15'h1EA8] =  8'hF4;
		ram[15'h1EA9] =  8'hB5;
		ram[15'h1EAA] =  8'h56;
		ram[15'h1EAB] =  8'hB3;
		ram[15'h1EAC] =  8'hC4;
		ram[15'h1EAD] =  8'h23;
		ram[15'h1EAE] =  8'hCF;
		ram[15'h1EAF] =  8'hBA;
		ram[15'h1EB0] =  8'h95;
		ram[15'h1EB1] =  8'h99;
		ram[15'h1EB2] =  8'hB8;
		ram[15'h1EB3] =  8'hBD;
		ram[15'h1EB4] =  8'hA5;
		ram[15'h1EB5] =  8'h0F;
		ram[15'h1EB6] =  8'h28;
		ram[15'h1EB7] =  8'h02;
		ram[15'h1EB8] =  8'hB8;
		ram[15'h1EB9] =  8'h9E;
		ram[15'h1EBA] =  8'h5F;
		ram[15'h1EBB] =  8'h05;
		ram[15'h1EBC] =  8'h88;
		ram[15'h1EBD] =  8'h08;
		ram[15'h1EBE] =  8'hC6;
		ram[15'h1EBF] =  8'h0C;
		ram[15'h1EC0] =  8'hD9;
		ram[15'h1EC1] =  8'hB2;
		ram[15'h1EC2] =  8'hB1;
		ram[15'h1EC3] =  8'h0B;
		ram[15'h1EC4] =  8'hE9;
		ram[15'h1EC5] =  8'h24;
		ram[15'h1EC6] =  8'h2F;
		ram[15'h1EC7] =  8'h6F;
		ram[15'h1EC8] =  8'h7C;
		ram[15'h1EC9] =  8'h87;
		ram[15'h1ECA] =  8'h58;
		ram[15'h1ECB] =  8'h68;
		ram[15'h1ECC] =  8'h4C;
		ram[15'h1ECD] =  8'h11;
		ram[15'h1ECE] =  8'hC1;
		ram[15'h1ECF] =  8'h61;
		ram[15'h1ED0] =  8'h1D;
		ram[15'h1ED1] =  8'hAB;
		ram[15'h1ED2] =  8'hB6;
		ram[15'h1ED3] =  8'h66;
		ram[15'h1ED4] =  8'h2D;
		ram[15'h1ED5] =  8'h3D;
		ram[15'h1ED6] =  8'h76;
		ram[15'h1ED7] =  8'hDC;
		ram[15'h1ED8] =  8'h41;
		ram[15'h1ED9] =  8'h90;
		ram[15'h1EDA] =  8'h01;
		ram[15'h1EDB] =  8'hDB;
		ram[15'h1EDC] =  8'h71;
		ram[15'h1EDD] =  8'h06;
		ram[15'h1EDE] =  8'h98;
		ram[15'h1EDF] =  8'hD2;
		ram[15'h1EE0] =  8'h20;
		ram[15'h1EE1] =  8'hBC;
		ram[15'h1EE2] =  8'hEF;
		ram[15'h1EE3] =  8'hD5;
		ram[15'h1EE4] =  8'h10;
		ram[15'h1EE5] =  8'h2A;
		ram[15'h1EE6] =  8'h71;
		ram[15'h1EE7] =  8'hB1;
		ram[15'h1EE8] =  8'h85;
		ram[15'h1EE9] =  8'h89;
		ram[15'h1EEA] =  8'h06;
		ram[15'h1EEB] =  8'hB6;
		ram[15'h1EEC] =  8'hB5;
		ram[15'h1EED] =  8'h1F;
		ram[15'h1EEE] =  8'h9F;
		ram[15'h1EEF] =  8'hBF;
		ram[15'h1EF0] =  8'hE4;
		ram[15'h1EF1] =  8'hA5;
		ram[15'h1EF2] =  8'hE8;
		ram[15'h1EF3] =  8'hB8;
		ram[15'h1EF4] =  8'hD4;
		ram[15'h1EF5] =  8'h33;
		ram[15'h1EF6] =  8'h78;
		ram[15'h1EF7] =  8'h07;
		ram[15'h1EF8] =  8'hC9;
		ram[15'h1EF9] =  8'hA2;
		ram[15'h1EFA] =  8'h0F;
		ram[15'h1EFB] =  8'h00;
		ram[15'h1EFC] =  8'hF9;
		ram[15'h1EFD] =  8'h34;
		ram[15'h1EFE] =  8'h96;
		ram[15'h1EFF] =  8'h09;
		ram[15'h1F00] =  8'hA8;
		ram[15'h1F01] =  8'h8E;
		ram[15'h1F02] =  8'hE1;
		ram[15'h1F03] =  8'h0E;
		ram[15'h1F04] =  8'h98;
		ram[15'h1F05] =  8'h18;
		ram[15'h1F06] =  8'h7F;
		ram[15'h1F07] =  8'h6A;
		ram[15'h1F08] =  8'h0D;
		ram[15'h1F09] =  8'hBB;
		ram[15'h1F0A] =  8'h08;
		ram[15'h1F0B] =  8'h6D;
		ram[15'h1F0C] =  8'h3D;
		ram[15'h1F0D] =  8'h2D;
		ram[15'h1F0E] =  8'h91;
		ram[15'h1F0F] =  8'h64;
		ram[15'h1F10] =  8'h6C;
		ram[15'h1F11] =  8'h97;
		ram[15'h1F12] =  8'hE6;
		ram[15'h1F13] =  8'h63;
		ram[15'h1F14] =  8'h5C;
		ram[15'h1F15] =  8'h01;
		ram[15'h1F16] =  8'h6B;
		ram[15'h1F17] =  8'h6B;
		ram[15'h1F18] =  8'h51;
		ram[15'h1F19] =  8'hF4;
		ram[15'h1F1A] =  8'h1C;
		ram[15'h1F1B] =  8'h6C;
		ram[15'h1F1C] =  8'h61;
		ram[15'h1F1D] =  8'h62;
		ram[15'h1F1E] =  8'h85;
		ram[15'h1F1F] =  8'h65;
		ram[15'h1F20] =  8'h30;
		ram[15'h1F21] =  8'hD8;
		ram[15'h1F22] =  8'hF2;
		ram[15'h1F23] =  8'h62;
		ram[15'h1F24] =  8'h00;
		ram[15'h1F25] =  8'h4E;
		ram[15'h1F26] =  8'h6C;
		ram[15'h1F27] =  8'h06;
		ram[15'h1F28] =  8'h95;
		ram[15'h1F29] =  8'hED;
		ram[15'h1F2A] =  8'h1B;
		ram[15'h1F2B] =  8'h01;
		ram[15'h1F2C] =  8'hA5;
		ram[15'h1F2D] =  8'h7B;
		ram[15'h1F2E] =  8'h82;
		ram[15'h1F2F] =  8'h08;
		ram[15'h1F30] =  8'hF4;
		ram[15'h1F31] =  8'hC1;
		ram[15'h1F32] =  8'hF5;
		ram[15'h1F33] =  8'h0F;
		ram[15'h1F34] =  8'hC4;
		ram[15'h1F35] =  8'h57;
		ram[15'h1F36] =  8'h65;
		ram[15'h1F37] =  8'hB0;
		ram[15'h1F38] =  8'hD9;
		ram[15'h1F39] =  8'hC6;
		ram[15'h1F3A] =  8'h12;
		ram[15'h1F3B] =  8'hB7;
		ram[15'h1F3C] =  8'hE9;
		ram[15'h1F3D] =  8'h50;
		ram[15'h1F3E] =  8'h8B;
		ram[15'h1F3F] =  8'hBE;
		ram[15'h1F40] =  8'hB8;
		ram[15'h1F41] =  8'hEA;
		ram[15'h1F42] =  8'hFC;
		ram[15'h1F43] =  8'hB9;
		ram[15'h1F44] =  8'h88;
		ram[15'h1F45] =  8'h7C;
		ram[15'h1F46] =  8'h62;
		ram[15'h1F47] =  8'hDD;
		ram[15'h1F48] =  8'h1D;
		ram[15'h1F49] =  8'hDF;
		ram[15'h1F4A] =  8'h15;
		ram[15'h1F4B] =  8'hDA;
		ram[15'h1F4C] =  8'h2D;
		ram[15'h1F4D] =  8'h49;
		ram[15'h1F4E] =  8'h8C;
		ram[15'h1F4F] =  8'hD3;
		ram[15'h1F50] =  8'h7C;
		ram[15'h1F51] =  8'hF3;
		ram[15'h1F52] =  8'hFB;
		ram[15'h1F53] =  8'hD4;
		ram[15'h1F54] =  8'h4C;
		ram[15'h1F55] =  8'h65;
		ram[15'h1F56] =  8'h4D;
		ram[15'h1F57] =  8'hB2;
		ram[15'h1F58] =  8'h61;
		ram[15'h1F59] =  8'h58;
		ram[15'h1F5A] =  8'h3A;
		ram[15'h1F5B] =  8'hB5;
		ram[15'h1F5C] =  8'h51;
		ram[15'h1F5D] =  8'hCE;
		ram[15'h1F5E] =  8'hA3;
		ram[15'h1F5F] =  8'hBC;
		ram[15'h1F60] =  8'h00;
		ram[15'h1F61] =  8'h74;
		ram[15'h1F62] =  8'hD4;
		ram[15'h1F63] =  8'hBB;
		ram[15'h1F64] =  8'h30;
		ram[15'h1F65] =  8'hE2;
		ram[15'h1F66] =  8'h4A;
		ram[15'h1F67] =  8'hDF;
		ram[15'h1F68] =  8'hA5;
		ram[15'h1F69] =  8'h41;
		ram[15'h1F6A] =  8'h3D;
		ram[15'h1F6B] =  8'hD8;
		ram[15'h1F6C] =  8'h95;
		ram[15'h1F6D] =  8'hD7;
		ram[15'h1F6E] =  8'hA4;
		ram[15'h1F6F] =  8'hD1;
		ram[15'h1F70] =  8'hC4;
		ram[15'h1F71] =  8'h6D;
		ram[15'h1F72] =  8'hD3;
		ram[15'h1F73] =  8'hD6;
		ram[15'h1F74] =  8'hF4;
		ram[15'h1F75] =  8'hFB;
		ram[15'h1F76] =  8'h43;
		ram[15'h1F77] =  8'h69;
		ram[15'h1F78] =  8'hE9;
		ram[15'h1F79] =  8'h6A;
		ram[15'h1F7A] =  8'h34;
		ram[15'h1F7B] =  8'h6E;
		ram[15'h1F7C] =  8'hD9;
		ram[15'h1F7D] =  8'hFC;
		ram[15'h1F7E] =  8'hAD;
		ram[15'h1F7F] =  8'h67;
		ram[15'h1F80] =  8'h88;
		ram[15'h1F81] =  8'h46;
		ram[15'h1F82] =  8'hDA;
		ram[15'h1F83] =  8'h60;
		ram[15'h1F84] =  8'hB8;
		ram[15'h1F85] =  8'hD0;
		ram[15'h1F86] =  8'h44;
		ram[15'h1F87] =  8'h04;
		ram[15'h1F88] =  8'h2D;
		ram[15'h1F89] =  8'h73;
		ram[15'h1F8A] =  8'h33;
		ram[15'h1F8B] =  8'h03;
		ram[15'h1F8C] =  8'h1D;
		ram[15'h1F8D] =  8'hE5;
		ram[15'h1F8E] =  8'hAA;
		ram[15'h1F8F] =  8'h0A;
		ram[15'h1F90] =  8'h4C;
		ram[15'h1F91] =  8'h5F;
		ram[15'h1F92] =  8'hDD;
		ram[15'h1F93] =  8'h0D;
		ram[15'h1F94] =  8'h7C;
		ram[15'h1F95] =  8'hC9;
		ram[15'h1F96] =  8'h50;
		ram[15'h1F97] =  8'h05;
		ram[15'h1F98] =  8'h71;
		ram[15'h1F99] =  8'h3C;
		ram[15'h1F9A] =  8'h27;
		ram[15'h1F9B] =  8'h02;
		ram[15'h1F9C] =  8'h41;
		ram[15'h1F9D] =  8'hAA;
		ram[15'h1F9E] =  8'hBE;
		ram[15'h1F9F] =  8'h0B;
		ram[15'h1FA0] =  8'h10;
		ram[15'h1FA1] =  8'h10;
		ram[15'h1FA2] =  8'hC9;
		ram[15'h1FA3] =  8'h0C;
		ram[15'h1FA4] =  8'h20;
		ram[15'h1FA5] =  8'h86;
		ram[15'h1FA6] =  8'h57;
		ram[15'h1FA7] =  8'h68;
		ram[15'h1FA8] =  8'hB5;
		ram[15'h1FA9] =  8'h25;
		ram[15'h1FAA] =  8'h20;
		ram[15'h1FAB] =  8'h6F;
		ram[15'h1FAC] =  8'h85;
		ram[15'h1FAD] =  8'hB3;
		ram[15'h1FAE] =  8'hB9;
		ram[15'h1FAF] =  8'h66;
		ram[15'h1FB0] =  8'hD4;
		ram[15'h1FB1] =  8'h09;
		ram[15'h1FB2] =  8'hCE;
		ram[15'h1FB3] =  8'h61;
		ram[15'h1FB4] =  8'hE4;
		ram[15'h1FB5] =  8'h9F;
		ram[15'h1FB6] =  8'h5E;
		ram[15'h1FB7] =  8'hDE;
		ram[15'h1FB8] =  8'hF9;
		ram[15'h1FB9] =  8'h0E;
		ram[15'h1FBA] =  8'h29;
		ram[15'h1FBB] =  8'hD9;
		ram[15'h1FBC] =  8'hC9;
		ram[15'h1FBD] =  8'h98;
		ram[15'h1FBE] =  8'hB0;
		ram[15'h1FBF] =  8'hD0;
		ram[15'h1FC0] =  8'h98;
		ram[15'h1FC1] =  8'h22;
		ram[15'h1FC2] =  8'hC7;
		ram[15'h1FC3] =  8'hD7;
		ram[15'h1FC4] =  8'hA8;
		ram[15'h1FC5] =  8'hB4;
		ram[15'h1FC6] =  8'h59;
		ram[15'h1FC7] =  8'hB3;
		ram[15'h1FC8] =  8'h3D;
		ram[15'h1FC9] =  8'h17;
		ram[15'h1FCA] =  8'h2E;
		ram[15'h1FCB] =  8'hB4;
		ram[15'h1FCC] =  8'h0D;
		ram[15'h1FCD] =  8'h81;
		ram[15'h1FCE] =  8'hB7;
		ram[15'h1FCF] =  8'hBD;
		ram[15'h1FD0] =  8'h5C;
		ram[15'h1FD1] =  8'h3B;
		ram[15'h1FD2] =  8'hC0;
		ram[15'h1FD3] =  8'hBA;
		ram[15'h1FD4] =  8'h6C;
		ram[15'h1FD5] =  8'hAD;
		ram[15'h1FD6] =  8'hED;
		ram[15'h1FD7] =  8'hB8;
		ram[15'h1FD8] =  8'h83;
		ram[15'h1FD9] =  8'h20;
		ram[15'h1FDA] =  8'h9A;
		ram[15'h1FDB] =  8'hBF;
		ram[15'h1FDC] =  8'hB3;
		ram[15'h1FDD] =  8'hB6;
		ram[15'h1FDE] =  8'h03;
		ram[15'h1FDF] =  8'hB6;
		ram[15'h1FE0] =  8'hE2;
		ram[15'h1FE1] =  8'h0C;
		ram[15'h1FE2] =  8'h74;
		ram[15'h1FE3] =  8'hB1;
		ram[15'h1FE4] =  8'hD2;
		ram[15'h1FE5] =  8'h9A;
		ram[15'h1FE6] =  8'hEA;
		ram[15'h1FE7] =  8'hD5;
		ram[15'h1FE8] =  8'h47;
		ram[15'h1FE9] =  8'h39;
		ram[15'h1FEA] =  8'h9D;
		ram[15'h1FEB] =  8'hD2;
		ram[15'h1FEC] =  8'h77;
		ram[15'h1FED] =  8'hAF;
		ram[15'h1FEE] =  8'h04;
		ram[15'h1FEF] =  8'hDB;
		ram[15'h1FF0] =  8'h26;
		ram[15'h1FF1] =  8'h15;
		ram[15'h1FF2] =  8'h73;
		ram[15'h1FF3] =  8'hDC;
		ram[15'h1FF4] =  8'h16;
		ram[15'h1FF5] =  8'h83;
		ram[15'h1FF6] =  8'hE3;
		ram[15'h1FF7] =  8'h63;
		ram[15'h1FF8] =  8'h0B;
		ram[15'h1FF9] =  8'h12;
		ram[15'h1FFA] =  8'h94;
		ram[15'h1FFB] =  8'h64;
		ram[15'h1FFC] =  8'h3B;
		ram[15'h1FFD] =  8'h84;
		ram[15'h1FFE] =  8'h0D;
		ram[15'h1FFF] =  8'h6D;
		ram[15'h2000] =  8'h6A;
		ram[15'h2001] =  8'h3E;
		ram[15'h2002] =  8'h7A;
		ram[15'h2003] =  8'h6A;
		ram[15'h2004] =  8'h5A;
		ram[15'h2005] =  8'hA8;
		ram[15'h2006] =  8'hE4;
		ram[15'h2007] =  8'h0E;
		ram[15'h2008] =  8'hCF;
		ram[15'h2009] =  8'h0B;
		ram[15'h200A] =  8'h93;
		ram[15'h200B] =  8'h09;
		ram[15'h200C] =  8'hFF;
		ram[15'h200D] =  8'h9D;
		ram[15'h200E] =  8'h0A;
		ram[15'h200F] =  8'h00;
		ram[15'h2010] =  8'hAE;
		ram[15'h2011] =  8'h27;
		ram[15'h2012] =  8'h7D;
		ram[15'h2013] =  8'h07;
		ram[15'h2014] =  8'h9E;
		ram[15'h2015] =  8'hB1;
		ram[15'h2016] =  8'hF0;
		ram[15'h2017] =  8'h0F;
		ram[15'h2018] =  8'h93;
		ram[15'h2019] =  8'h44;
		ram[15'h201A] =  8'h87;
		ram[15'h201B] =  8'h08;
		ram[15'h201C] =  8'hA3;
		ram[15'h201D] =  8'hD2;
		ram[15'h201E] =  8'h1E;
		ram[15'h201F] =  8'h01;
		ram[15'h2020] =  8'hF2;
		ram[15'h2021] =  8'h68;
		ram[15'h2022] =  8'h69;
		ram[15'h2023] =  8'h06;
		ram[15'h2024] =  8'hC2;
		ram[15'h2025] =  8'hFE;
		ram[15'h2026] =  8'hF7;
		ram[15'h2027] =  8'h62;
		ram[15'h2028] =  8'h57;
		ram[15'h2029] =  8'h5D;
		ram[15'h202A] =  8'h80;
		ram[15'h202B] =  8'h65;
		ram[15'h202C] =  8'h67;
		ram[15'h202D] =  8'hCB;
		ram[15'h202E] =  8'h19;
		ram[15'h202F] =  8'h6C;
		ram[15'h2030] =  8'h36;
		ram[15'h2031] =  8'h71;
		ram[15'h2032] =  8'h6E;
		ram[15'h2033] =  8'h6B;
		ram[15'h2034] =  8'h06;
		ram[15'h2035] =  8'hE7;
		ram[15'h2036] =  8'hFE;
		ram[15'h2037] =  8'hD4;
		ram[15'h2038] =  8'h1B;
		ram[15'h2039] =  8'h76;
		ram[15'h203A] =  8'h89;
		ram[15'h203B] =  8'hD3;
		ram[15'h203C] =  8'h2B;
		ram[15'h203D] =  8'hE0;
		ram[15'h203E] =  8'h10;
		ram[15'h203F] =  8'hDA;
		ram[15'h2040] =  8'h7A;
		ram[15'h2041] =  8'h5A;
		ram[15'h2042] =  8'h67;
		ram[15'h2043] =  8'hDD;
		ram[15'h2044] =  8'h4A;
		ram[15'h2045] =  8'hCC;
		ram[15'h2046] =  8'hF9;
		ram[15'h2047] =  8'hB9;
		ram[15'h2048] =  8'hDF;
		ram[15'h2049] =  8'h6F;
		ram[15'h204A] =  8'h8E;
		ram[15'h204B] =  8'hBE;
		ram[15'h204C] =  8'hEF;
		ram[15'h204D] =  8'hF9;
		ram[15'h204E] =  8'h17;
		ram[15'h204F] =  8'hB7;
		ram[15'h2050] =  8'hBE;
		ram[15'h2051] =  8'h43;
		ram[15'h2052] =  8'h60;
		ram[15'h2053] =  8'hB0;
		ram[15'h2054] =  8'h8E;
		ram[15'h2055] =  8'hD5;
		ram[15'h2056] =  8'hD6;
		ram[15'h2057] =  8'hD6;
		ram[15'h2058] =  8'hA3;
		ram[15'h2059] =  8'hE8;
		ram[15'h205A] =  8'hA1;
		ram[15'h205B] =  8'hD1;
		ram[15'h205C] =  8'h93;
		ram[15'h205D] =  8'h7E;
		ram[15'h205E] =  8'h38;
		ram[15'h205F] =  8'hD8;
		ram[15'h2060] =  8'hC2;
		ram[15'h2061] =  8'hC4;
		ram[15'h2062] =  8'h4F;
		ram[15'h2063] =  8'hDF;
		ram[15'h2064] =  8'hF2;
		ram[15'h2065] =  8'h52;
		ram[15'h2066] =  8'hD1;
		ram[15'h2067] =  8'hBB;
		ram[15'h2068] =  8'h67;
		ram[15'h2069] =  8'hF1;
		ram[15'h206A] =  8'hA6;
		ram[15'h206B] =  8'hBC;
		ram[15'h206C] =  8'h57;
		ram[15'h206D] =  8'h67;
		ram[15'h206E] =  8'h3F;
		ram[15'h206F] =  8'hB5;
		ram[15'h2070] =  8'h06;
		ram[15'h2071] =  8'hDD;
		ram[15'h2072] =  8'h48;
		ram[15'h2073] =  8'hB2;
		ram[15'h2074] =  8'h36;
		ram[15'h2075] =  8'h4B;
		ram[15'h2076] =  8'hD8;
		ram[15'h2077] =  8'h0D;
		ram[15'h2078] =  8'h2B;
		ram[15'h2079] =  8'hDA;
		ram[15'h207A] =  8'hAF;
		ram[15'h207B] =  8'h0A;
		ram[15'h207C] =  8'h1B;
		ram[15'h207D] =  8'h4C;
		ram[15'h207E] =  8'h36;
		ram[15'h207F] =  8'h03;
		ram[15'h2080] =  8'h4A;
		ram[15'h2081] =  8'hF6;
		ram[15'h2082] =  8'h41;
		ram[15'h2083] =  8'h04;
		ram[15'h2084] =  8'h7A;
		ram[15'h2085] =  8'h60;
		ram[15'h2086] =  8'hDF;
		ram[15'h2087] =  8'h60;
		ram[15'h2088] =  8'hEF;
		ram[15'h2089] =  8'hC3;
		ram[15'h208A] =  8'hA8;
		ram[15'h208B] =  8'h67;
		ram[15'h208C] =  8'hDF;
		ram[15'h208D] =  8'h55;
		ram[15'h208E] =  8'h31;
		ram[15'h208F] =  8'h6E;
		ram[15'h2090] =  8'h8E;
		ram[15'h2091] =  8'hEF;
		ram[15'h2092] =  8'h46;
		ram[15'h2093] =  8'h69;
		ram[15'h2094] =  8'hBE;
		ram[15'h2095] =  8'h79;
		ram[15'h2096] =  8'hCB;
		ram[15'h2097] =  8'h61;
		ram[15'h2098] =  8'hB3;
		ram[15'h2099] =  8'h8C;
		ram[15'h209A] =  8'hBC;
		ram[15'h209B] =  8'h66;
		ram[15'h209C] =  8'h83;
		ram[15'h209D] =  8'h1A;
		ram[15'h209E] =  8'h25;
		ram[15'h209F] =  8'h6F;
		ram[15'h20A0] =  8'hD2;
		ram[15'h20A1] =  8'hA0;
		ram[15'h20A2] =  8'h52;
		ram[15'h20A3] =  8'h68;
		ram[15'h20A4] =  8'hE2;
		ram[15'h20A5] =  8'h36;
		ram[15'h20A6] =  8'hCC;
		ram[15'h20A7] =  8'h0C;
		ram[15'h20A8] =  8'h77;
		ram[15'h20A9] =  8'h95;
		ram[15'h20AA] =  8'hBB;
		ram[15'h20AB] =  8'h0B;
		ram[15'h20AC] =  8'h47;
		ram[15'h20AD] =  8'h03;
		ram[15'h20AE] =  8'h22;
		ram[15'h20AF] =  8'h02;
		ram[15'h20B0] =  8'h16;
		ram[15'h20B1] =  8'hB9;
		ram[15'h20B2] =  8'h55;
		ram[15'h20B3] =  8'h05;
		ram[15'h20B4] =  8'h26;
		ram[15'h20B5] =  8'h2F;
		ram[15'h20B6] =  8'hC5;
		ram[15'h20B7] =  8'hBA;
		ram[15'h20B8] =  8'h3B;
		ram[15'h20B9] =  8'hBE;
		ram[15'h20BA] =  8'hB2;
		ram[15'h20BB] =  8'hBD;
		ram[15'h20BC] =  8'h0B;
		ram[15'h20BD] =  8'h28;
		ram[15'h20BE] =  8'h2B;
		ram[15'h20BF] =  8'hB4;
		ram[15'h20C0] =  8'h5A;
		ram[15'h20C1] =  8'h92;
		ram[15'h20C2] =  8'h5C;
		ram[15'h20C3] =  8'hB3;
		ram[15'h20C4] =  8'h6A;
		ram[15'h20C5] =  8'h04;
		ram[15'h20C6] =  8'hC2;
		ram[15'h20C7] =  8'hD7;
		ram[15'h20C8] =  8'hFF;
		ram[15'h20C9] =  8'hA7;
		ram[15'h20CA] =  8'hB5;
		ram[15'h20CB] =  8'hD0;
		ram[15'h20CC] =  8'hCF;
		ram[15'h20CD] =  8'h31;
		ram[15'h20CE] =  8'h2C;
		ram[15'h20CF] =  8'hD9;
		ram[15'h20D0] =  8'h9E;
		ram[15'h20D1] =  8'h8B;
		ram[15'h20D2] =  8'h5B;
		ram[15'h20D3] =  8'hDE;
		ram[15'h20D4] =  8'hAE;
		ram[15'h20D5] =  8'h1D;
		ram[15'h20D6] =  8'h9B;
		ram[15'h20D7] =  8'h64;
		ram[15'h20D8] =  8'hC2;
		ram[15'h20D9] =  8'hB0;
		ram[15'h20DA] =  8'hEC;
		ram[15'h20DB] =  8'h63;
		ram[15'h20DC] =  8'hF2;
		ram[15'h20DD] =  8'h26;
		ram[15'h20DE] =  8'h75;
		ram[15'h20DF] =  8'h6A;
		ram[15'h20E0] =  8'hA3;
		ram[15'h20E1] =  8'h9C;
		ram[15'h20E2] =  8'h02;
		ram[15'h20E3] =  8'h6D;
		ram[15'h20E4] =  8'h93;
		ram[15'h20E5] =  8'h0A;
		ram[15'h20E6] =  8'h9C;
		ram[15'h20E7] =  8'h09;
		ram[15'h20E8] =  8'h06;
		ram[15'h20E9] =  8'hA9;
		ram[15'h20EA] =  8'hEB;
		ram[15'h20EB] =  8'h0E;
		ram[15'h20EC] =  8'h36;
		ram[15'h20ED] =  8'h3F;
		ram[15'h20EE] =  8'h72;
		ram[15'h20EF] =  8'h07;
		ram[15'h20F0] =  8'h67;
		ram[15'h20F1] =  8'h85;
		ram[15'h20F2] =  8'h05;
		ram[15'h20F3] =  8'h00;
		ram[15'h20F4] =  8'h57;
		ram[15'h20F5] =  8'h13;
		ram[15'h20F6] =  8'h95;
		ram[15'h20F7] =  8'hBF;
		ram[15'h20F8] =  8'h4A;
		ram[15'h20F9] =  8'h82;
		ram[15'h20FA] =  8'hE2;
		ram[15'h20FB] =  8'hB8;
		ram[15'h20FC] =  8'h7A;
		ram[15'h20FD] =  8'h14;
		ram[15'h20FE] =  8'h7B;
		ram[15'h20FF] =  8'hB1;
		ram[15'h2100] =  8'h2B;
		ram[15'h2101] =  8'hAE;
		ram[15'h2102] =  8'h0C;
		ram[15'h2103] =  8'hB6;
		ram[15'h2104] =  8'h1B;
		ram[15'h2105] =  8'h38;
		ram[15'h2106] =  8'h92;
		ram[15'h2107] =  8'hD2;
		ram[15'h2108] =  8'h8E;
		ram[15'h2109] =  8'h9B;
		ram[15'h210A] =  8'hE5;
		ram[15'h210B] =  8'hD5;
		ram[15'h210C] =  8'hBE;
		ram[15'h210D] =  8'h0D;
		ram[15'h210E] =  8'h7C;
		ram[15'h210F] =  8'hDC;
		ram[15'h2110] =  8'hEF;
		ram[15'h2111] =  8'hB7;
		ram[15'h2112] =  8'h0B;
		ram[15'h2113] =  8'hDB;
		ram[15'h2114] =  8'hDF;
		ram[15'h2115] =  8'h21;
		ram[15'h2116] =  8'h86;
		ram[15'h2117] =  8'hD3;
		ram[15'h2118] =  8'hD2;
		ram[15'h2119] =  8'hD4;
		ram[15'h211A] =  8'hF1;
		ram[15'h211B] =  8'hD4;
		ram[15'h211C] =  8'hE2;
		ram[15'h211D] =  8'h42;
		ram[15'h211E] =  8'h68;
		ram[15'h211F] =  8'hDD;
		ram[15'h2120] =  8'hB3;
		ram[15'h2121] =  8'hF8;
		ram[15'h2122] =  8'h1F;
		ram[15'h2123] =  8'hDA;
		ram[15'h2124] =  8'h83;
		ram[15'h2125] =  8'h6E;
		ram[15'h2126] =  8'h81;
		ram[15'h2127] =  8'hBE;
		ram[15'h2128] =  8'h16;
		ram[15'h2129] =  8'hCD;
		ram[15'h212A] =  8'hF6;
		ram[15'h212B] =  8'hB9;
		ram[15'h212C] =  8'h26;
		ram[15'h212D] =  8'h5B;
		ram[15'h212E] =  8'h6F;
		ram[15'h212F] =  8'hB0;
		ram[15'h2130] =  8'h77;
		ram[15'h2131] =  8'hE1;
		ram[15'h2132] =  8'h18;
		ram[15'h2133] =  8'hB7;
		ram[15'h2134] =  8'h47;
		ram[15'h2135] =  8'h77;
		ram[15'h2136] =  8'h88;
		ram[15'h2137] =  8'h08;
		ram[15'h2138] =  8'h5A;
		ram[15'h2139] =  8'hE6;
		ram[15'h213A] =  8'hFF;
		ram[15'h213B] =  8'h0F;
		ram[15'h213C] =  8'h6A;
		ram[15'h213D] =  8'h70;
		ram[15'h213E] =  8'h66;
		ram[15'h213F] =  8'h06;
		ram[15'h2140] =  8'h3B;
		ram[15'h2141] =  8'hCA;
		ram[15'h2142] =  8'h11;
		ram[15'h2143] =  8'h01;
		ram[15'h2144] =  8'h0B;
		ram[15'h2145] =  8'h5C;
		ram[15'h2146] =  8'h8F;
		ram[15'h2147] =  8'h65;
		ram[15'h2148] =  8'h9E;
		ram[15'h2149] =  8'hFF;
		ram[15'h214A] =  8'hF8;
		ram[15'h214B] =  8'h62;
		ram[15'h214C] =  8'hAE;
		ram[15'h214D] =  8'h69;
		ram[15'h214E] =  8'h61;
		ram[15'h214F] =  8'h6B;
		ram[15'h2150] =  8'hFF;
		ram[15'h2151] =  8'hD3;
		ram[15'h2152] =  8'h16;
		ram[15'h2153] =  8'h6C;
		ram[15'h2154] =  8'hCF;
		ram[15'h2155] =  8'h45;
		ram[15'h2156] =  8'hA0;
		ram[15'h2157] =  8'h0A;
		ram[15'h2158] =  8'hE2;
		ram[15'h2159] =  8'h78;
		ram[15'h215A] =  8'hD7;
		ram[15'h215B] =  8'h0D;
		ram[15'h215C] =  8'hD2;
		ram[15'h215D] =  8'hEE;
		ram[15'h215E] =  8'h4E;
		ram[15'h215F] =  8'h04;
		ram[15'h2160] =  8'h83;
		ram[15'h2161] =  8'h54;
		ram[15'h2162] =  8'h39;
		ram[15'h2163] =  8'h03;
		ram[15'h2164] =  8'hB3;
		ram[15'h2165] =  8'hC2;
		ram[15'h2166] =  8'hA7;
		ram[15'h2167] =  8'h67;
		ram[15'h2168] =  8'h26;
		ram[15'h2169] =  8'h61;
		ram[15'h216A] =  8'hD0;
		ram[15'h216B] =  8'h60;
		ram[15'h216C] =  8'h16;
		ram[15'h216D] =  8'hF7;
		ram[15'h216E] =  8'h49;
		ram[15'h216F] =  8'h69;
		ram[15'h2170] =  8'h47;
		ram[15'h2171] =  8'h4D;
		ram[15'h2172] =  8'h3E;
		ram[15'h2173] =  8'h6E;
		ram[15'h2174] =  8'h77;
		ram[15'h2175] =  8'hDB;
		ram[15'h2176] =  8'hAE;
		ram[15'h2177] =  8'hD1;
		ram[15'h2178] =  8'h6A;
		ram[15'h2179] =  8'h4A;
		ram[15'h217A] =  8'hD9;
		ram[15'h217B] =  8'hD6;
		ram[15'h217C] =  8'h5A;
		ram[15'h217D] =  8'hDC;
		ram[15'h217E] =  8'h40;
		ram[15'h217F] =  8'hDF;
		ram[15'h2180] =  8'h0B;
		ram[15'h2181] =  8'h66;
		ram[15'h2182] =  8'h37;
		ram[15'h2183] =  8'hD8;
		ram[15'h2184] =  8'h3B;
		ram[15'h2185] =  8'hF0;
		ram[15'h2186] =  8'hA9;
		ram[15'h2187] =  8'hBC;
		ram[15'h2188] =  8'hAE;
		ram[15'h2189] =  8'h53;
		ram[15'h218A] =  8'hDE;
		ram[15'h218B] =  8'hBB;
		ram[15'h218C] =  8'h9E;
		ram[15'h218D] =  8'hC5;
		ram[15'h218E] =  8'h47;
		ram[15'h218F] =  8'hB2;
		ram[15'h2190] =  8'hCF;
		ram[15'h2191] =  8'h7F;
		ram[15'h2192] =  8'h30;
		ram[15'h2193] =  8'hB5;
		ram[15'h2194] =  8'hFF;
		ram[15'h2195] =  8'hE9;
		ram[15'h2196] =  8'hBD;
		ram[15'h2197] =  8'hBD;
		ram[15'h2198] =  8'hF2;
		ram[15'h2199] =  8'h1C;
		ram[15'h219A] =  8'hCA;
		ram[15'h219B] =  8'hBA;
		ram[15'h219C] =  8'hC2;
		ram[15'h219D] =  8'h8A;
		ram[15'h219E] =  8'h53;
		ram[15'h219F] =  8'hB3;
		ram[15'h21A0] =  8'h93;
		ram[15'h21A1] =  8'h30;
		ram[15'h21A2] =  8'h24;
		ram[15'h21A3] =  8'hB4;
		ram[15'h21A4] =  8'hA3;
		ram[15'h21A5] =  8'hA6;
		ram[15'h21A6] =  8'hBA;
		ram[15'h21A7] =  8'hD0;
		ram[15'h21A8] =  8'h36;
		ram[15'h21A9] =  8'h05;
		ram[15'h21AA] =  8'hCD;
		ram[15'h21AB] =  8'hD7;
		ram[15'h21AC] =  8'h06;
		ram[15'h21AD] =  8'h93;
		ram[15'h21AE] =  8'h54;
		ram[15'h21AF] =  8'hDE;
		ram[15'h21B0] =  8'h57;
		ram[15'h21B1] =  8'h29;
		ram[15'h21B2] =  8'h23;
		ram[15'h21B3] =  8'hD9;
		ram[15'h21B4] =  8'h67;
		ram[15'h21B5] =  8'hBF;
		ram[15'h21B6] =  8'hB3;
		ram[15'h21B7] =  8'h66;
		ram[15'h21B8] =  8'h7A;
		ram[15'h21B9] =  8'h2E;
		ram[15'h21BA] =  8'hC4;
		ram[15'h21BB] =  8'h61;
		ram[15'h21BC] =  8'h4A;
		ram[15'h21BD] =  8'hB8;
		ram[15'h21BE] =  8'h5D;
		ram[15'h21BF] =  8'h68;
		ram[15'h21C0] =  8'h1B;
		ram[15'h21C1] =  8'h02;
		ram[15'h21C2] =  8'h2A;
		ram[15'h21C3] =  8'h6F;
		ram[15'h21C4] =  8'h2B;
		ram[15'h21C5] =  8'h94;
		ram[15'h21C6] =  8'hB4;
		ram[15'h21C7] =  8'h0B;
		ram[15'h21C8] =  8'hBE;
		ram[15'h21C9] =  8'h37;
		ram[15'h21CA] =  8'hC3;
		ram[15'h21CB] =  8'h0C;
		ram[15'h21CC] =  8'h8E;
		ram[15'h21CD] =  8'hA1;
		ram[15'h21CE] =  8'h5A;
		ram[15'h21CF] =  8'h05;
		ram[15'h21D0] =  8'hDF;
		ram[15'h21D1] =  8'h1B;
		ram[15'h21D2] =  8'h2D;
		ram[15'h21D3] =  8'h02;
		ram[15'h21D4] =  8'hEF;
		ram[15'h21D5] =  8'h8D;

		
end

endmodule 