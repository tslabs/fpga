module top
(
	input wire DCLK,
	input wire DATA0
);
	
	sfl	sfl
	(
		.noe_in	(1'b0)
	);
	
endmodule
