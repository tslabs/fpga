`timescale 1ns / 1ps

module ssram(
	input	wire		CLK,
	
	input	wire [14:0]	ADDR, //16kb
	input	wire [7:0]	DI,
	output	wire [7:0]	DO,
	input	wire		OE,
	input	wire		WE
); 	   

reg [7:0]	ram [0:32*1024-1];

always @ (negedge CLK)
if (WE)		 	
begin
	ram[ADDR] = DI;
	//$display("MEM WRITE ADDR=%h VAL=%h", ADDR, DI);
end
	
assign #1 DO = ram[ADDR];

integer i;

initial
begin	
		for(i=0;i<32*1024;i=i+1)
			ram[i] = 0;
	
		
		
		
		
		ram[15'h0] = 8'hF3;
		ram[15'h1] = 8'h18;
		ram[15'h2] = 8'h37;
		ram[15'h3] = 8'h00;
		ram[15'h4] = 8'h00;
		ram[15'h5] = 8'h00;
		ram[15'h6] = 8'h00;
		ram[15'h7] = 8'h00;
		ram[15'h8] = 8'h00;
		ram[15'h9] = 8'h00;
		ram[15'hA] = 8'h00;
		ram[15'hB] = 8'h00;
		ram[15'hC] = 8'h00;
		ram[15'hD] = 8'h00;
		ram[15'hE] = 8'h00;
		ram[15'hF] = 8'h00;
		ram[15'h10] = 8'hD3;
		ram[15'h11] = 8'hFF;
		ram[15'h12] = 8'hC9;
		ram[15'h13] = 8'h00;
		ram[15'h14] = 8'h00;
		ram[15'h15] = 8'h00;
		ram[15'h16] = 8'h00;
		ram[15'h17] = 8'h00;
		ram[15'h18] = 8'hC9;
		ram[15'h19] = 8'h00;
		ram[15'h1A] = 8'h00;
		ram[15'h1B] = 8'h00;
		ram[15'h1C] = 8'h00;
		ram[15'h1D] = 8'h00;
		ram[15'h1E] = 8'h00;
		ram[15'h1F] = 8'h00;
		ram[15'h20] = 8'hED;
		ram[15'h21] = 8'h4D;
		ram[15'h22] = 8'h00;
		ram[15'h23] = 8'h00;
		ram[15'h24] = 8'h00;
		ram[15'h25] = 8'h00;
		ram[15'h26] = 8'h00;
		ram[15'h27] = 8'h00;
		ram[15'h28] = 8'hED;
		ram[15'h29] = 8'h45;
		ram[15'h2A] = 8'h00;
		ram[15'h2B] = 8'h00;
		ram[15'h2C] = 8'h00;
		ram[15'h2D] = 8'h00;
		ram[15'h2E] = 8'h00;
		ram[15'h2F] = 8'h00;
		ram[15'h30] = 8'h00;
		ram[15'h31] = 8'h00;
		ram[15'h32] = 8'h00;
		ram[15'h33] = 8'h00;
		ram[15'h34] = 8'h00;
		ram[15'h35] = 8'h00;
		ram[15'h36] = 8'h00;
		ram[15'h37] = 8'h00;
		ram[15'h38] = 8'hED;
		ram[15'h39] = 8'h4D;
		ram[15'h3A] = 8'h21;
		ram[15'h3B] = 8'hEC;
		ram[15'h3C] = 8'h0C;
		ram[15'h3D] = 8'hF9;
		ram[15'h3E] = 8'h00;
		ram[15'h3F] = 8'h00;
		ram[15'h40] = 8'h21;
		ram[15'h41] = 8'h00;
		ram[15'h42] = 8'h00;
		ram[15'h43] = 8'h11;
		ram[15'h44] = 8'h00;
		ram[15'h45] = 8'h00;
		ram[15'h46] = 8'h01;
		ram[15'h47] = 8'h00;
		ram[15'h48] = 8'h00;
		ram[15'h49] = 8'hC5;
		ram[15'h4A] = 8'hF1;
		ram[15'h4B] = 8'hDD;
		ram[15'h4C] = 8'h21;
		ram[15'h4D] = 8'h00;
		ram[15'h4E] = 8'h00;
		ram[15'h4F] = 8'hFD;
		ram[15'h50] = 8'h21;
		ram[15'h51] = 8'h00;
		ram[15'h52] = 8'h00;
		ram[15'h53] = 8'hE5;
		ram[15'h54] = 8'hD5;
		ram[15'h55] = 8'hC5;
		ram[15'h56] = 8'hD9;
		ram[15'h57] = 8'hC1;
		ram[15'h58] = 8'hD1;
		ram[15'h59] = 8'hE1;
		ram[15'h5A] = 8'hD9;
		ram[15'h5B] = 8'hFB;
		ram[15'h5C] = 8'hCD;
		ram[15'h5D] = 8'hA8;
		ram[15'h5E] = 8'h00;
		ram[15'h5F] = 8'hCD;
		ram[15'h60] = 8'h4E;
		ram[15'h61] = 8'h01;
		ram[15'h62] = 8'hCD;
		ram[15'h63] = 8'h81;
		ram[15'h64] = 8'h01;
		ram[15'h65] = 8'hCD;
		ram[15'h66] = 8'hAA;
		ram[15'h67] = 8'h01;
		ram[15'h68] = 8'hCD;
		ram[15'h69] = 8'h34;
		ram[15'h6A] = 8'h02;
		ram[15'h6B] = 8'hCD;
		ram[15'h6C] = 8'h55;
		ram[15'h6D] = 8'h02;
		ram[15'h6E] = 8'hCD;
		ram[15'h6F] = 8'hC3;
		ram[15'h70] = 8'h02;
		ram[15'h71] = 8'hCD;
		ram[15'h72] = 8'hF3;
		ram[15'h73] = 8'h02;
		ram[15'h74] = 8'hCD;
		ram[15'h75] = 8'hC2;
		ram[15'h76] = 8'h03;
		ram[15'h77] = 8'hCD;
		ram[15'h78] = 8'h6C;
		ram[15'h79] = 8'h05;
		ram[15'h7A] = 8'hCD;
		ram[15'h7B] = 8'h82;
		ram[15'h7C] = 8'h05;
		ram[15'h7D] = 8'hCD;
		ram[15'h7E] = 8'h87;
		ram[15'h7F] = 8'h05;
		ram[15'h80] = 8'hCD;
		ram[15'h81] = 8'h5A;
		ram[15'h82] = 8'h06;
		ram[15'h83] = 8'hCD;
		ram[15'h84] = 8'h7B;
		ram[15'h85] = 8'h07;
		ram[15'h86] = 8'hCD;
		ram[15'h87] = 8'h6E;
		ram[15'h88] = 8'h0A;
		ram[15'h89] = 8'hCD;
		ram[15'h8A] = 8'h09;
		ram[15'h8B] = 8'h0B;
		ram[15'h8C] = 8'hCD;
		ram[15'h8D] = 8'hDC;
		ram[15'h8E] = 8'h0B;
		ram[15'h8F] = 8'h76;
		ram[15'h90] = 8'h18;
		ram[15'h91] = 8'hFD;
		ram[15'h92] = 8'h00;
		ram[15'h93] = 8'h00;
		ram[15'h94] = 8'h00;
		ram[15'h95] = 8'h00;
		ram[15'h96] = 8'h00;
		ram[15'h97] = 8'h00;
		ram[15'h98] = 8'h00;
		ram[15'h99] = 8'h00;
		ram[15'h9A] = 8'h00;
		ram[15'h9B] = 8'h00;
		ram[15'h9C] = 8'h00;
		ram[15'h9D] = 8'h00;
		ram[15'h9E] = 8'h00;
		ram[15'h9F] = 8'h00;
		ram[15'hA0] = 8'h00;
		ram[15'hA1] = 8'h00;
		ram[15'hA2] = 8'h00;
		ram[15'hA3] = 8'h00;
		ram[15'hA4] = 8'h00;
		ram[15'hA5] = 8'h00;
		ram[15'hA6] = 8'h00;
		ram[15'hA7] = 8'h00;
		ram[15'hA8] = 8'h3E;
		ram[15'hA9] = 8'h01;
		ram[15'hAA] = 8'hD3;
		ram[15'hAB] = 8'h01;
		ram[15'hAC] = 8'h3E;
		ram[15'hAD] = 8'h07;
		ram[15'hAE] = 8'h77;
		ram[15'hAF] = 8'h01;
		ram[15'hB0] = 8'h02;
		ram[15'hB1] = 8'h01;
		ram[15'hB2] = 8'h11;
		ram[15'hB3] = 8'h04;
		ram[15'hB4] = 8'h03;
		ram[15'hB5] = 8'h21;
		ram[15'hB6] = 8'h06;
		ram[15'hB7] = 8'h05;
		ram[15'hB8] = 8'h78;
		ram[15'hB9] = 8'h79;
		ram[15'hBA] = 8'h7A;
		ram[15'hBB] = 8'h7B;
		ram[15'hBC] = 8'h7C;
		ram[15'hBD] = 8'h7D;
		ram[15'hBE] = 8'h21;
		ram[15'hBF] = 8'h92;
		ram[15'hC0] = 8'h00;
		ram[15'hC1] = 8'h7E;
		ram[15'hC2] = 8'h7F;
		ram[15'hC3] = 8'h3E;
		ram[15'hC4] = 8'h07;
		ram[15'hC5] = 8'h40;
		ram[15'hC6] = 8'h41;
		ram[15'hC7] = 8'h42;
		ram[15'hC8] = 8'h43;
		ram[15'hC9] = 8'h44;
		ram[15'hCA] = 8'h45;
		ram[15'hCB] = 8'h21;
		ram[15'hCC] = 8'h92;
		ram[15'hCD] = 8'h00;
		ram[15'hCE] = 8'h46;
		ram[15'hCF] = 8'h47;
		ram[15'hD0] = 8'h06;
		ram[15'hD1] = 8'h01;
		ram[15'hD2] = 8'h48;
		ram[15'hD3] = 8'h49;
		ram[15'hD4] = 8'h4A;
		ram[15'hD5] = 8'h4B;
		ram[15'hD6] = 8'h4C;
		ram[15'hD7] = 8'h4D;
		ram[15'hD8] = 8'h21;
		ram[15'hD9] = 8'h92;
		ram[15'hDA] = 8'h00;
		ram[15'hDB] = 8'h4E;
		ram[15'hDC] = 8'h4F;
		ram[15'hDD] = 8'h0E;
		ram[15'hDE] = 8'h02;
		ram[15'hDF] = 8'h50;
		ram[15'hE0] = 8'h51;
		ram[15'hE1] = 8'h52;
		ram[15'hE2] = 8'h53;
		ram[15'hE3] = 8'h54;
		ram[15'hE4] = 8'h55;
		ram[15'hE5] = 8'h21;
		ram[15'hE6] = 8'h92;
		ram[15'hE7] = 8'h00;
		ram[15'hE8] = 8'h56;
		ram[15'hE9] = 8'h57;
		ram[15'hEA] = 8'h16;
		ram[15'hEB] = 8'h03;
		ram[15'hEC] = 8'h58;
		ram[15'hED] = 8'h59;
		ram[15'hEE] = 8'h5A;
		ram[15'hEF] = 8'h5B;
		ram[15'hF0] = 8'h5C;
		ram[15'hF1] = 8'h5D;
		ram[15'hF2] = 8'h21;
		ram[15'hF3] = 8'h92;
		ram[15'hF4] = 8'h00;
		ram[15'hF5] = 8'h5E;
		ram[15'hF6] = 8'h5F;
		ram[15'hF7] = 8'h1E;
		ram[15'hF8] = 8'h04;
		ram[15'hF9] = 8'h60;
		ram[15'hFA] = 8'h61;
		ram[15'hFB] = 8'h62;
		ram[15'hFC] = 8'h63;
		ram[15'hFD] = 8'h64;
		ram[15'hFE] = 8'h65;
		ram[15'hFF] = 8'h21;
		ram[15'h100] = 8'h92;
		ram[15'h101] = 8'h00;
		ram[15'h102] = 8'h66;
		ram[15'h103] = 8'h67;
		ram[15'h104] = 8'h26;
		ram[15'h105] = 8'h05;
		ram[15'h106] = 8'h68;
		ram[15'h107] = 8'h69;
		ram[15'h108] = 8'h6A;
		ram[15'h109] = 8'h6B;
		ram[15'h10A] = 8'h6C;
		ram[15'h10B] = 8'h6D;
		ram[15'h10C] = 8'h21;
		ram[15'h10D] = 8'h92;
		ram[15'h10E] = 8'h00;
		ram[15'h10F] = 8'h6E;
		ram[15'h110] = 8'h6F;
		ram[15'h111] = 8'h21;
		ram[15'h112] = 8'h92;
		ram[15'h113] = 8'h00;
		ram[15'h114] = 8'h70;
		ram[15'h115] = 8'h71;
		ram[15'h116] = 8'h72;
		ram[15'h117] = 8'h73;
		ram[15'h118] = 8'h74;
		ram[15'h119] = 8'h75;
		ram[15'h11A] = 8'h77;
		ram[15'h11B] = 8'hDD;
		ram[15'h11C] = 8'h21;
		ram[15'h11D] = 8'h92;
		ram[15'h11E] = 8'h00;
		ram[15'h11F] = 8'hDD;
		ram[15'h120] = 8'h70;
		ram[15'h121] = 8'h00;
		ram[15'h122] = 8'hDD;
		ram[15'h123] = 8'h71;
		ram[15'h124] = 8'h01;
		ram[15'h125] = 8'hDD;
		ram[15'h126] = 8'h72;
		ram[15'h127] = 8'h02;
		ram[15'h128] = 8'hDD;
		ram[15'h129] = 8'h73;
		ram[15'h12A] = 8'h03;
		ram[15'h12B] = 8'hDD;
		ram[15'h12C] = 8'h74;
		ram[15'h12D] = 8'h00;
		ram[15'h12E] = 8'hDD;
		ram[15'h12F] = 8'h75;
		ram[15'h130] = 8'h01;
		ram[15'h131] = 8'hDD;
		ram[15'h132] = 8'h77;
		ram[15'h133] = 8'h02;
		ram[15'h134] = 8'hFD;
		ram[15'h135] = 8'h21;
		ram[15'h136] = 8'h92;
		ram[15'h137] = 8'h00;
		ram[15'h138] = 8'hFD;
		ram[15'h139] = 8'h46;
		ram[15'h13A] = 8'h00;
		ram[15'h13B] = 8'hFD;
		ram[15'h13C] = 8'h4E;
		ram[15'h13D] = 8'h01;
		ram[15'h13E] = 8'hFD;
		ram[15'h13F] = 8'h56;
		ram[15'h140] = 8'h02;
		ram[15'h141] = 8'hFD;
		ram[15'h142] = 8'h5E;
		ram[15'h143] = 8'h03;
		ram[15'h144] = 8'hFD;
		ram[15'h145] = 8'h66;
		ram[15'h146] = 8'h00;
		ram[15'h147] = 8'hFD;
		ram[15'h148] = 8'h6E;
		ram[15'h149] = 8'h01;
		ram[15'h14A] = 8'hFD;
		ram[15'h14B] = 8'h7E;
		ram[15'h14C] = 8'h02;
		ram[15'h14D] = 8'hC9;
		ram[15'h14E] = 8'h3E;
		ram[15'h14F] = 8'h02;
		ram[15'h150] = 8'hD3;
		ram[15'h151] = 8'h01;
		ram[15'h152] = 8'h3E;
		ram[15'h153] = 8'h01;
		ram[15'h154] = 8'h32;
		ram[15'h155] = 8'h92;
		ram[15'h156] = 8'h00;
		ram[15'h157] = 8'h06;
		ram[15'h158] = 8'h02;
		ram[15'h159] = 8'h78;
		ram[15'h15A] = 8'h32;
		ram[15'h15B] = 8'h92;
		ram[15'h15C] = 8'h00;
		ram[15'h15D] = 8'h0E;
		ram[15'h15E] = 8'h03;
		ram[15'h15F] = 8'h79;
		ram[15'h160] = 8'h32;
		ram[15'h161] = 8'h92;
		ram[15'h162] = 8'h00;
		ram[15'h163] = 8'h16;
		ram[15'h164] = 8'h04;
		ram[15'h165] = 8'h7A;
		ram[15'h166] = 8'h32;
		ram[15'h167] = 8'h92;
		ram[15'h168] = 8'h00;
		ram[15'h169] = 8'h1E;
		ram[15'h16A] = 8'h05;
		ram[15'h16B] = 8'h7B;
		ram[15'h16C] = 8'h32;
		ram[15'h16D] = 8'h92;
		ram[15'h16E] = 8'h00;
		ram[15'h16F] = 8'h26;
		ram[15'h170] = 8'h04;
		ram[15'h171] = 8'h32;
		ram[15'h172] = 8'h92;
		ram[15'h173] = 8'h00;
		ram[15'h174] = 8'h7C;
		ram[15'h175] = 8'h2E;
		ram[15'h176] = 8'h05;
		ram[15'h177] = 8'h7D;
		ram[15'h178] = 8'h32;
		ram[15'h179] = 8'h92;
		ram[15'h17A] = 8'h00;
		ram[15'h17B] = 8'h21;
		ram[15'h17C] = 8'h92;
		ram[15'h17D] = 8'h00;
		ram[15'h17E] = 8'h36;
		ram[15'h17F] = 8'h06;
		ram[15'h180] = 8'hC9;
		ram[15'h181] = 8'h3E;
		ram[15'h182] = 8'h03;
		ram[15'h183] = 8'hD3;
		ram[15'h184] = 8'h01;
		ram[15'h185] = 8'h01;
		ram[15'h186] = 8'h02;
		ram[15'h187] = 8'h01;
		ram[15'h188] = 8'hED;
		ram[15'h189] = 8'h43;
		ram[15'h18A] = 8'h96;
		ram[15'h18B] = 8'h00;
		ram[15'h18C] = 8'h11;
		ram[15'h18D] = 8'h04;
		ram[15'h18E] = 8'h03;
		ram[15'h18F] = 8'hED;
		ram[15'h190] = 8'h53;
		ram[15'h191] = 8'h96;
		ram[15'h192] = 8'h00;
		ram[15'h193] = 8'h21;
		ram[15'h194] = 8'h06;
		ram[15'h195] = 8'h05;
		ram[15'h196] = 8'h22;
		ram[15'h197] = 8'h96;
		ram[15'h198] = 8'h00;
		ram[15'h199] = 8'hDD;
		ram[15'h19A] = 8'h21;
		ram[15'h19B] = 8'h08;
		ram[15'h19C] = 8'h07;
		ram[15'h19D] = 8'hDD;
		ram[15'h19E] = 8'h22;
		ram[15'h19F] = 8'h96;
		ram[15'h1A0] = 8'h00;
		ram[15'h1A1] = 8'hFD;
		ram[15'h1A2] = 8'h21;
		ram[15'h1A3] = 8'h0A;
		ram[15'h1A4] = 8'h09;
		ram[15'h1A5] = 8'hFD;
		ram[15'h1A6] = 8'h22;
		ram[15'h1A7] = 8'h96;
		ram[15'h1A8] = 8'h00;
		ram[15'h1A9] = 8'hC9;
		ram[15'h1AA] = 8'h3E;
		ram[15'h1AB] = 8'h04;
		ram[15'h1AC] = 8'hD3;
		ram[15'h1AD] = 8'h01;
		ram[15'h1AE] = 8'h01;
		ram[15'h1AF] = 8'h02;
		ram[15'h1B0] = 8'h01;
		ram[15'h1B1] = 8'h11;
		ram[15'h1B2] = 8'h04;
		ram[15'h1B3] = 8'h03;
		ram[15'h1B4] = 8'h21;
		ram[15'h1B5] = 8'h06;
		ram[15'h1B6] = 8'h05;
		ram[15'h1B7] = 8'h3E;
		ram[15'h1B8] = 8'h07;
		ram[15'h1B9] = 8'hDD;
		ram[15'h1BA] = 8'h21;
		ram[15'h1BB] = 8'h92;
		ram[15'h1BC] = 8'h00;
		ram[15'h1BD] = 8'hFD;
		ram[15'h1BE] = 8'h21;
		ram[15'h1BF] = 8'h92;
		ram[15'h1C0] = 8'h00;
		ram[15'h1C1] = 8'hDD;
		ram[15'h1C2] = 8'h77;
		ram[15'h1C3] = 8'h00;
		ram[15'h1C4] = 8'hDD;
		ram[15'h1C5] = 8'h70;
		ram[15'h1C6] = 8'h01;
		ram[15'h1C7] = 8'hDD;
		ram[15'h1C8] = 8'h71;
		ram[15'h1C9] = 8'h02;
		ram[15'h1CA] = 8'hDD;
		ram[15'h1CB] = 8'h72;
		ram[15'h1CC] = 8'h03;
		ram[15'h1CD] = 8'hDD;
		ram[15'h1CE] = 8'h73;
		ram[15'h1CF] = 8'h00;
		ram[15'h1D0] = 8'hDD;
		ram[15'h1D1] = 8'h74;
		ram[15'h1D2] = 8'h01;
		ram[15'h1D3] = 8'hDD;
		ram[15'h1D4] = 8'h75;
		ram[15'h1D5] = 8'h02;
		ram[15'h1D6] = 8'hFD;
		ram[15'h1D7] = 8'h21;
		ram[15'h1D8] = 8'h92;
		ram[15'h1D9] = 8'h00;
		ram[15'h1DA] = 8'hFD;
		ram[15'h1DB] = 8'h77;
		ram[15'h1DC] = 8'h03;
		ram[15'h1DD] = 8'hFD;
		ram[15'h1DE] = 8'h70;
		ram[15'h1DF] = 8'h00;
		ram[15'h1E0] = 8'hFD;
		ram[15'h1E1] = 8'h71;
		ram[15'h1E2] = 8'h01;
		ram[15'h1E3] = 8'hFD;
		ram[15'h1E4] = 8'h72;
		ram[15'h1E5] = 8'h02;
		ram[15'h1E6] = 8'hFD;
		ram[15'h1E7] = 8'h73;
		ram[15'h1E8] = 8'h03;
		ram[15'h1E9] = 8'hFD;
		ram[15'h1EA] = 8'h74;
		ram[15'h1EB] = 8'h00;
		ram[15'h1EC] = 8'hFD;
		ram[15'h1ED] = 8'h75;
		ram[15'h1EE] = 8'h01;
		ram[15'h1EF] = 8'h21;
		ram[15'h1F0] = 8'h92;
		ram[15'h1F1] = 8'h00;
		ram[15'h1F2] = 8'h36;
		ram[15'h1F3] = 8'h01;
		ram[15'h1F4] = 8'h23;
		ram[15'h1F5] = 8'h36;
		ram[15'h1F6] = 8'h02;
		ram[15'h1F7] = 8'h23;
		ram[15'h1F8] = 8'h36;
		ram[15'h1F9] = 8'h03;
		ram[15'h1FA] = 8'h23;
		ram[15'h1FB] = 8'h36;
		ram[15'h1FC] = 8'h04;
		ram[15'h1FD] = 8'hDD;
		ram[15'h1FE] = 8'h7E;
		ram[15'h1FF] = 8'h00;
		ram[15'h200] = 8'hDD;
		ram[15'h201] = 8'h46;
		ram[15'h202] = 8'h01;
		ram[15'h203] = 8'hDD;
		ram[15'h204] = 8'h4E;
		ram[15'h205] = 8'h02;
		ram[15'h206] = 8'hDD;
		ram[15'h207] = 8'h56;
		ram[15'h208] = 8'h03;
		ram[15'h209] = 8'hDD;
		ram[15'h20A] = 8'h5E;
		ram[15'h20B] = 8'h00;
		ram[15'h20C] = 8'hDD;
		ram[15'h20D] = 8'h66;
		ram[15'h20E] = 8'h01;
		ram[15'h20F] = 8'hDD;
		ram[15'h210] = 8'h6E;
		ram[15'h211] = 8'h02;
		ram[15'h212] = 8'hFD;
		ram[15'h213] = 8'h7E;
		ram[15'h214] = 8'h03;
		ram[15'h215] = 8'hFD;
		ram[15'h216] = 8'h46;
		ram[15'h217] = 8'h00;
		ram[15'h218] = 8'hFD;
		ram[15'h219] = 8'h4E;
		ram[15'h21A] = 8'h01;
		ram[15'h21B] = 8'hFD;
		ram[15'h21C] = 8'h56;
		ram[15'h21D] = 8'h02;
		ram[15'h21E] = 8'hFD;
		ram[15'h21F] = 8'h5E;
		ram[15'h220] = 8'h03;
		ram[15'h221] = 8'hFD;
		ram[15'h222] = 8'h66;
		ram[15'h223] = 8'h00;
		ram[15'h224] = 8'hFD;
		ram[15'h225] = 8'h6E;
		ram[15'h226] = 8'h01;
		ram[15'h227] = 8'hDD;
		ram[15'h228] = 8'h36;
		ram[15'h229] = 8'h01;
		ram[15'h22A] = 8'h10;
		ram[15'h22B] = 8'hFD;
		ram[15'h22C] = 8'h36;
		ram[15'h22D] = 8'h02;
		ram[15'h22E] = 8'h11;
		ram[15'h22F] = 8'hDD;
		ram[15'h230] = 8'h36;
		ram[15'h231] = 8'h03;
		ram[15'h232] = 8'h13;
		ram[15'h233] = 8'hC9;
		ram[15'h234] = 8'h3E;
		ram[15'h235] = 8'h05;
		ram[15'h236] = 8'hD3;
		ram[15'h237] = 8'h01;
		ram[15'h238] = 8'h01;
		ram[15'h239] = 8'h92;
		ram[15'h23A] = 8'h00;
		ram[15'h23B] = 8'h11;
		ram[15'h23C] = 8'h93;
		ram[15'h23D] = 8'h00;
		ram[15'h23E] = 8'h3E;
		ram[15'h23F] = 8'h20;
		ram[15'h240] = 8'h02;
		ram[15'h241] = 8'h3E;
		ram[15'h242] = 8'h21;
		ram[15'h243] = 8'h12;
		ram[15'h244] = 8'h0A;
		ram[15'h245] = 8'h1A;
		ram[15'h246] = 8'h32;
		ram[15'h247] = 8'h92;
		ram[15'h248] = 8'h00;
		ram[15'h249] = 8'h3A;
		ram[15'h24A] = 8'h92;
		ram[15'h24B] = 8'h00;
		ram[15'h24C] = 8'hED;
		ram[15'h24D] = 8'h57;
		ram[15'h24E] = 8'hED;
		ram[15'h24F] = 8'h47;
		ram[15'h250] = 8'hED;
		ram[15'h251] = 8'h5F;
		ram[15'h252] = 8'hED;
		ram[15'h253] = 8'h4F;
		ram[15'h254] = 8'hC9;
		ram[15'h255] = 8'h3E;
		ram[15'h256] = 8'h06;
		ram[15'h257] = 8'hD3;
		ram[15'h258] = 8'h01;
		ram[15'h259] = 8'h01;
		ram[15'h25A] = 8'h02;
		ram[15'h25B] = 8'h01;
		ram[15'h25C] = 8'hED;
		ram[15'h25D] = 8'h43;
		ram[15'h25E] = 8'h96;
		ram[15'h25F] = 8'h00;
		ram[15'h260] = 8'hED;
		ram[15'h261] = 8'h4B;
		ram[15'h262] = 8'h96;
		ram[15'h263] = 8'h00;
		ram[15'h264] = 8'h11;
		ram[15'h265] = 8'h04;
		ram[15'h266] = 8'h03;
		ram[15'h267] = 8'hED;
		ram[15'h268] = 8'h53;
		ram[15'h269] = 8'h96;
		ram[15'h26A] = 8'h00;
		ram[15'h26B] = 8'hED;
		ram[15'h26C] = 8'h5B;
		ram[15'h26D] = 8'h96;
		ram[15'h26E] = 8'h00;
		ram[15'h26F] = 8'h21;
		ram[15'h270] = 8'h06;
		ram[15'h271] = 8'h05;
		ram[15'h272] = 8'h22;
		ram[15'h273] = 8'h96;
		ram[15'h274] = 8'h00;
		ram[15'h275] = 8'h2A;
		ram[15'h276] = 8'h96;
		ram[15'h277] = 8'h00;
		ram[15'h278] = 8'hF3;
		ram[15'h279] = 8'hED;
		ram[15'h27A] = 8'h73;
		ram[15'h27B] = 8'h96;
		ram[15'h27C] = 8'h00;
		ram[15'h27D] = 8'hCD;
		ram[15'h27E] = 8'h80;
		ram[15'h27F] = 8'h02;
		ram[15'h280] = 8'hE1;
		ram[15'h281] = 8'h31;
		ram[15'h282] = 8'h00;
		ram[15'h283] = 8'h00;
		ram[15'h284] = 8'hF9;
		ram[15'h285] = 8'hE5;
		ram[15'h286] = 8'hDD;
		ram[15'h287] = 8'hE1;
		ram[15'h288] = 8'hDD;
		ram[15'h289] = 8'hF9;
		ram[15'h28A] = 8'hE5;
		ram[15'h28B] = 8'hFD;
		ram[15'h28C] = 8'hE1;
		ram[15'h28D] = 8'hFD;
		ram[15'h28E] = 8'hF9;
		ram[15'h28F] = 8'hED;
		ram[15'h290] = 8'h7B;
		ram[15'h291] = 8'h96;
		ram[15'h292] = 8'h00;
		ram[15'h293] = 8'hFB;
		ram[15'h294] = 8'hDD;
		ram[15'h295] = 8'h21;
		ram[15'h296] = 8'h08;
		ram[15'h297] = 8'h07;
		ram[15'h298] = 8'hDD;
		ram[15'h299] = 8'h22;
		ram[15'h29A] = 8'h96;
		ram[15'h29B] = 8'h00;
		ram[15'h29C] = 8'hDD;
		ram[15'h29D] = 8'h2A;
		ram[15'h29E] = 8'h96;
		ram[15'h29F] = 8'h00;
		ram[15'h2A0] = 8'hFD;
		ram[15'h2A1] = 8'h21;
		ram[15'h2A2] = 8'h0A;
		ram[15'h2A3] = 8'h09;
		ram[15'h2A4] = 8'hFD;
		ram[15'h2A5] = 8'h22;
		ram[15'h2A6] = 8'h96;
		ram[15'h2A7] = 8'h00;
		ram[15'h2A8] = 8'hFD;
		ram[15'h2A9] = 8'h2A;
		ram[15'h2AA] = 8'h96;
		ram[15'h2AB] = 8'h00;
		ram[15'h2AC] = 8'h2A;
		ram[15'h2AD] = 8'h96;
		ram[15'h2AE] = 8'h00;
		ram[15'h2AF] = 8'hC5;
		ram[15'h2B0] = 8'hD5;
		ram[15'h2B1] = 8'hE5;
		ram[15'h2B2] = 8'hF5;
		ram[15'h2B3] = 8'hDD;
		ram[15'h2B4] = 8'hE5;
		ram[15'h2B5] = 8'hFD;
		ram[15'h2B6] = 8'hE5;
		ram[15'h2B7] = 8'hF3;
		ram[15'h2B8] = 8'h00;
		ram[15'h2B9] = 8'hFB;
		ram[15'h2BA] = 8'hFD;
		ram[15'h2BB] = 8'hE1;
		ram[15'h2BC] = 8'hDD;
		ram[15'h2BD] = 8'hE1;
		ram[15'h2BE] = 8'hF1;
		ram[15'h2BF] = 8'hE1;
		ram[15'h2C0] = 8'hD1;
		ram[15'h2C1] = 8'hC1;
		ram[15'h2C2] = 8'hC9;
		ram[15'h2C3] = 8'h3E;
		ram[15'h2C4] = 8'h07;
		ram[15'h2C5] = 8'hD3;
		ram[15'h2C6] = 8'h01;
		ram[15'h2C7] = 8'h11;
		ram[15'h2C8] = 8'h02;
		ram[15'h2C9] = 8'h01;
		ram[15'h2CA] = 8'h21;
		ram[15'h2CB] = 8'h04;
		ram[15'h2CC] = 8'h03;
		ram[15'h2CD] = 8'hEB;
		ram[15'h2CE] = 8'h21;
		ram[15'h2CF] = 8'h20;
		ram[15'h2D0] = 8'h10;
		ram[15'h2D1] = 8'hE5;
		ram[15'h2D2] = 8'h21;
		ram[15'h2D3] = 8'h40;
		ram[15'h2D4] = 8'h30;
		ram[15'h2D5] = 8'hE5;
		ram[15'h2D6] = 8'hF1;
		ram[15'h2D7] = 8'h08;
		ram[15'h2D8] = 8'hF1;
		ram[15'h2D9] = 8'h08;
		ram[15'h2DA] = 8'h21;
		ram[15'h2DB] = 8'h60;
		ram[15'h2DC] = 8'h50;
		ram[15'h2DD] = 8'hE5;
		ram[15'h2DE] = 8'h21;
		ram[15'h2DF] = 8'h02;
		ram[15'h2E0] = 8'h01;
		ram[15'h2E1] = 8'hE3;
		ram[15'h2E2] = 8'h22;
		ram[15'h2E3] = 8'h96;
		ram[15'h2E4] = 8'h00;
		ram[15'h2E5] = 8'hDD;
		ram[15'h2E6] = 8'hE3;
		ram[15'h2E7] = 8'hDD;
		ram[15'h2E8] = 8'h22;
		ram[15'h2E9] = 8'h96;
		ram[15'h2EA] = 8'h00;
		ram[15'h2EB] = 8'hFD;
		ram[15'h2EC] = 8'hE3;
		ram[15'h2ED] = 8'hFD;
		ram[15'h2EE] = 8'h22;
		ram[15'h2EF] = 8'h96;
		ram[15'h2F0] = 8'h00;
		ram[15'h2F1] = 8'hE1;
		ram[15'h2F2] = 8'hC9;
		ram[15'h2F3] = 8'h3E;
		ram[15'h2F4] = 8'h08;
		ram[15'h2F5] = 8'hD3;
		ram[15'h2F6] = 8'h01;
		ram[15'h2F7] = 8'h21;
		ram[15'h2F8] = 8'h98;
		ram[15'h2F9] = 8'h00;
		ram[15'h2FA] = 8'h54;
		ram[15'h2FB] = 8'h5D;
		ram[15'h2FC] = 8'h13;
		ram[15'h2FD] = 8'h36;
		ram[15'h2FE] = 8'hAA;
		ram[15'h2FF] = 8'h01;
		ram[15'h300] = 8'h0F;
		ram[15'h301] = 8'h00;
		ram[15'h302] = 8'hED;
		ram[15'h303] = 8'hB0;
		ram[15'h304] = 8'h22;
		ram[15'h305] = 8'h96;
		ram[15'h306] = 8'h00;
		ram[15'h307] = 8'hED;
		ram[15'h308] = 8'h53;
		ram[15'h309] = 8'h96;
		ram[15'h30A] = 8'h00;
		ram[15'h30B] = 8'hED;
		ram[15'h30C] = 8'h43;
		ram[15'h30D] = 8'h96;
		ram[15'h30E] = 8'h00;
		ram[15'h30F] = 8'h21;
		ram[15'h310] = 8'hA7;
		ram[15'h311] = 8'h00;
		ram[15'h312] = 8'h54;
		ram[15'h313] = 8'h5D;
		ram[15'h314] = 8'h1B;
		ram[15'h315] = 8'h01;
		ram[15'h316] = 8'h0F;
		ram[15'h317] = 8'h00;
		ram[15'h318] = 8'h36;
		ram[15'h319] = 8'h55;
		ram[15'h31A] = 8'hED;
		ram[15'h31B] = 8'hB8;
		ram[15'h31C] = 8'h22;
		ram[15'h31D] = 8'h96;
		ram[15'h31E] = 8'h00;
		ram[15'h31F] = 8'hED;
		ram[15'h320] = 8'h53;
		ram[15'h321] = 8'h96;
		ram[15'h322] = 8'h00;
		ram[15'h323] = 8'hED;
		ram[15'h324] = 8'h43;
		ram[15'h325] = 8'h96;
		ram[15'h326] = 8'h00;
		ram[15'h327] = 8'h21;
		ram[15'h328] = 8'h98;
		ram[15'h329] = 8'h00;
		ram[15'h32A] = 8'h11;
		ram[15'h32B] = 8'h99;
		ram[15'h32C] = 8'h00;
		ram[15'h32D] = 8'h01;
		ram[15'h32E] = 8'h0F;
		ram[15'h32F] = 8'h00;
		ram[15'h330] = 8'h36;
		ram[15'h331] = 8'h0F;
		ram[15'h332] = 8'hED;
		ram[15'h333] = 8'hA0;
		ram[15'h334] = 8'hED;
		ram[15'h335] = 8'hA0;
		ram[15'h336] = 8'hED;
		ram[15'h337] = 8'hA0;
		ram[15'h338] = 8'hED;
		ram[15'h339] = 8'hA0;
		ram[15'h33A] = 8'h22;
		ram[15'h33B] = 8'h96;
		ram[15'h33C] = 8'h00;
		ram[15'h33D] = 8'hED;
		ram[15'h33E] = 8'h53;
		ram[15'h33F] = 8'h96;
		ram[15'h340] = 8'h00;
		ram[15'h341] = 8'hED;
		ram[15'h342] = 8'h43;
		ram[15'h343] = 8'h96;
		ram[15'h344] = 8'h00;
		ram[15'h345] = 8'h21;
		ram[15'h346] = 8'hA7;
		ram[15'h347] = 8'h00;
		ram[15'h348] = 8'h11;
		ram[15'h349] = 8'hA6;
		ram[15'h34A] = 8'h00;
		ram[15'h34B] = 8'h01;
		ram[15'h34C] = 8'h0F;
		ram[15'h34D] = 8'h00;
		ram[15'h34E] = 8'h36;
		ram[15'h34F] = 8'hF0;
		ram[15'h350] = 8'hED;
		ram[15'h351] = 8'hA8;
		ram[15'h352] = 8'hED;
		ram[15'h353] = 8'hA8;
		ram[15'h354] = 8'hED;
		ram[15'h355] = 8'hA8;
		ram[15'h356] = 8'hED;
		ram[15'h357] = 8'hA8;
		ram[15'h358] = 8'h22;
		ram[15'h359] = 8'h96;
		ram[15'h35A] = 8'h00;
		ram[15'h35B] = 8'hED;
		ram[15'h35C] = 8'h53;
		ram[15'h35D] = 8'h96;
		ram[15'h35E] = 8'h00;
		ram[15'h35F] = 8'hED;
		ram[15'h360] = 8'h43;
		ram[15'h361] = 8'h96;
		ram[15'h362] = 8'h00;
		ram[15'h363] = 8'h21;
		ram[15'h364] = 8'h98;
		ram[15'h365] = 8'h00;
		ram[15'h366] = 8'h01;
		ram[15'h367] = 8'h0F;
		ram[15'h368] = 8'h00;
		ram[15'h369] = 8'h3E;
		ram[15'h36A] = 8'h0F;
		ram[15'h36B] = 8'hED;
		ram[15'h36C] = 8'hA1;
		ram[15'h36D] = 8'hED;
		ram[15'h36E] = 8'hA1;
		ram[15'h36F] = 8'hED;
		ram[15'h370] = 8'hA1;
		ram[15'h371] = 8'hED;
		ram[15'h372] = 8'hA1;
		ram[15'h373] = 8'hF5;
		ram[15'h374] = 8'hED;
		ram[15'h375] = 8'hA1;
		ram[15'h376] = 8'hF5;
		ram[15'h377] = 8'h00;
		ram[15'h378] = 8'hF1;
		ram[15'h379] = 8'hF1;
		ram[15'h37A] = 8'hED;
		ram[15'h37B] = 8'h43;
		ram[15'h37C] = 8'h96;
		ram[15'h37D] = 8'h00;
		ram[15'h37E] = 8'h22;
		ram[15'h37F] = 8'h96;
		ram[15'h380] = 8'h00;
		ram[15'h381] = 8'h21;
		ram[15'h382] = 8'hA7;
		ram[15'h383] = 8'h00;
		ram[15'h384] = 8'h01;
		ram[15'h385] = 8'h0F;
		ram[15'h386] = 8'h00;
		ram[15'h387] = 8'h3E;
		ram[15'h388] = 8'hF0;
		ram[15'h389] = 8'hED;
		ram[15'h38A] = 8'hA9;
		ram[15'h38B] = 8'hED;
		ram[15'h38C] = 8'hA9;
		ram[15'h38D] = 8'hED;
		ram[15'h38E] = 8'hA9;
		ram[15'h38F] = 8'hED;
		ram[15'h390] = 8'hA9;
		ram[15'h391] = 8'hF5;
		ram[15'h392] = 8'hED;
		ram[15'h393] = 8'hA9;
		ram[15'h394] = 8'hF5;
		ram[15'h395] = 8'h00;
		ram[15'h396] = 8'hF1;
		ram[15'h397] = 8'hF1;
		ram[15'h398] = 8'hED;
		ram[15'h399] = 8'h43;
		ram[15'h39A] = 8'h96;
		ram[15'h39B] = 8'h00;
		ram[15'h39C] = 8'h22;
		ram[15'h39D] = 8'h96;
		ram[15'h39E] = 8'h00;
		ram[15'h39F] = 8'h21;
		ram[15'h3A0] = 8'h98;
		ram[15'h3A1] = 8'h00;
		ram[15'h3A2] = 8'h01;
		ram[15'h3A3] = 8'h05;
		ram[15'h3A4] = 8'h00;
		ram[15'h3A5] = 8'h3E;
		ram[15'h3A6] = 8'h0F;
		ram[15'h3A7] = 8'hED;
		ram[15'h3A8] = 8'hB1;
		ram[15'h3A9] = 8'hED;
		ram[15'h3AA] = 8'h43;
		ram[15'h3AB] = 8'h96;
		ram[15'h3AC] = 8'h00;
		ram[15'h3AD] = 8'h22;
		ram[15'h3AE] = 8'h96;
		ram[15'h3AF] = 8'h00;
		ram[15'h3B0] = 8'h21;
		ram[15'h3B1] = 8'hA7;
		ram[15'h3B2] = 8'h00;
		ram[15'h3B3] = 8'h01;
		ram[15'h3B4] = 8'h05;
		ram[15'h3B5] = 8'h00;
		ram[15'h3B6] = 8'h3E;
		ram[15'h3B7] = 8'hF0;
		ram[15'h3B8] = 8'hED;
		ram[15'h3B9] = 8'hB9;
		ram[15'h3BA] = 8'hED;
		ram[15'h3BB] = 8'h43;
		ram[15'h3BC] = 8'h96;
		ram[15'h3BD] = 8'h00;
		ram[15'h3BE] = 8'h22;
		ram[15'h3BF] = 8'h96;
		ram[15'h3C0] = 8'h00;
		ram[15'h3C1] = 8'hC9;
		ram[15'h3C2] = 8'h3E;
		ram[15'h3C3] = 8'h09;
		ram[15'h3C4] = 8'hD3;
		ram[15'h3C5] = 8'h01;
		ram[15'h3C6] = 8'hDD;
		ram[15'h3C7] = 8'h21;
		ram[15'h3C8] = 8'h93;
		ram[15'h3C9] = 8'h00;
		ram[15'h3CA] = 8'hFD;
		ram[15'h3CB] = 8'h21;
		ram[15'h3CC] = 8'h93;
		ram[15'h3CD] = 8'h00;
		ram[15'h3CE] = 8'hDD;
		ram[15'h3CF] = 8'h36;
		ram[15'h3D0] = 8'h00;
		ram[15'h3D1] = 8'h09;
		ram[15'h3D2] = 8'hFD;
		ram[15'h3D3] = 8'h36;
		ram[15'h3D4] = 8'h00;
		ram[15'h3D5] = 8'h0A;
		ram[15'h3D6] = 8'h3E;
		ram[15'h3D7] = 8'h07;
		ram[15'h3D8] = 8'h01;
		ram[15'h3D9] = 8'h02;
		ram[15'h3DA] = 8'h01;
		ram[15'h3DB] = 8'h11;
		ram[15'h3DC] = 8'h04;
		ram[15'h3DD] = 8'h03;
		ram[15'h3DE] = 8'h21;
		ram[15'h3DF] = 8'h06;
		ram[15'h3E0] = 8'h05;
		ram[15'h3E1] = 8'h87;
		ram[15'h3E2] = 8'h80;
		ram[15'h3E3] = 8'h81;
		ram[15'h3E4] = 8'h82;
		ram[15'h3E5] = 8'h83;
		ram[15'h3E6] = 8'h84;
		ram[15'h3E7] = 8'h85;
		ram[15'h3E8] = 8'h21;
		ram[15'h3E9] = 8'h92;
		ram[15'h3EA] = 8'h00;
		ram[15'h3EB] = 8'h36;
		ram[15'h3EC] = 8'h08;
		ram[15'h3ED] = 8'h86;
		ram[15'h3EE] = 8'hDD;
		ram[15'h3EF] = 8'h8E;
		ram[15'h3F0] = 8'h00;
		ram[15'h3F1] = 8'hFD;
		ram[15'h3F2] = 8'h8E;
		ram[15'h3F3] = 8'h01;
		ram[15'h3F4] = 8'hC6;
		ram[15'h3F5] = 8'h0B;
		ram[15'h3F6] = 8'h32;
		ram[15'h3F7] = 8'h92;
		ram[15'h3F8] = 8'h00;
		ram[15'h3F9] = 8'h3E;
		ram[15'h3FA] = 8'h07;
		ram[15'h3FB] = 8'h21;
		ram[15'h3FC] = 8'h06;
		ram[15'h3FD] = 8'h05;
		ram[15'h3FE] = 8'h8F;
		ram[15'h3FF] = 8'h88;
		ram[15'h400] = 8'h89;
		ram[15'h401] = 8'h8A;
		ram[15'h402] = 8'h8B;
		ram[15'h403] = 8'h8C;
		ram[15'h404] = 8'h8D;
		ram[15'h405] = 8'h21;
		ram[15'h406] = 8'h92;
		ram[15'h407] = 8'h00;
		ram[15'h408] = 8'h36;
		ram[15'h409] = 8'h08;
		ram[15'h40A] = 8'h8E;
		ram[15'h40B] = 8'hDD;
		ram[15'h40C] = 8'h8E;
		ram[15'h40D] = 8'h00;
		ram[15'h40E] = 8'hFD;
		ram[15'h40F] = 8'h8E;
		ram[15'h410] = 8'h01;
		ram[15'h411] = 8'hCE;
		ram[15'h412] = 8'h0B;
		ram[15'h413] = 8'h32;
		ram[15'h414] = 8'h92;
		ram[15'h415] = 8'h00;
		ram[15'h416] = 8'h3E;
		ram[15'h417] = 8'h07;
		ram[15'h418] = 8'h21;
		ram[15'h419] = 8'h06;
		ram[15'h41A] = 8'h05;
		ram[15'h41B] = 8'h97;
		ram[15'h41C] = 8'h97;
		ram[15'h41D] = 8'h97;
		ram[15'h41E] = 8'h90;
		ram[15'h41F] = 8'h97;
		ram[15'h420] = 8'h91;
		ram[15'h421] = 8'h97;
		ram[15'h422] = 8'h92;
		ram[15'h423] = 8'h97;
		ram[15'h424] = 8'h93;
		ram[15'h425] = 8'h97;
		ram[15'h426] = 8'h94;
		ram[15'h427] = 8'h97;
		ram[15'h428] = 8'h95;
		ram[15'h429] = 8'h21;
		ram[15'h42A] = 8'h92;
		ram[15'h42B] = 8'h00;
		ram[15'h42C] = 8'h36;
		ram[15'h42D] = 8'h08;
		ram[15'h42E] = 8'h97;
		ram[15'h42F] = 8'h96;
		ram[15'h430] = 8'h97;
		ram[15'h431] = 8'hDD;
		ram[15'h432] = 8'h96;
		ram[15'h433] = 8'h00;
		ram[15'h434] = 8'h97;
		ram[15'h435] = 8'hFD;
		ram[15'h436] = 8'h96;
		ram[15'h437] = 8'h01;
		ram[15'h438] = 8'h97;
		ram[15'h439] = 8'hD6;
		ram[15'h43A] = 8'h0B;
		ram[15'h43B] = 8'h32;
		ram[15'h43C] = 8'h92;
		ram[15'h43D] = 8'h00;
		ram[15'h43E] = 8'h3E;
		ram[15'h43F] = 8'h07;
		ram[15'h440] = 8'h21;
		ram[15'h441] = 8'h06;
		ram[15'h442] = 8'h05;
		ram[15'h443] = 8'h9F;
		ram[15'h444] = 8'h98;
		ram[15'h445] = 8'h99;
		ram[15'h446] = 8'h9A;
		ram[15'h447] = 8'h9B;
		ram[15'h448] = 8'h9C;
		ram[15'h449] = 8'h9D;
		ram[15'h44A] = 8'h21;
		ram[15'h44B] = 8'h92;
		ram[15'h44C] = 8'h00;
		ram[15'h44D] = 8'h36;
		ram[15'h44E] = 8'h08;
		ram[15'h44F] = 8'h9E;
		ram[15'h450] = 8'hDD;
		ram[15'h451] = 8'h9E;
		ram[15'h452] = 8'h00;
		ram[15'h453] = 8'hFD;
		ram[15'h454] = 8'h9E;
		ram[15'h455] = 8'h01;
		ram[15'h456] = 8'hDE;
		ram[15'h457] = 8'h0B;
		ram[15'h458] = 8'h32;
		ram[15'h459] = 8'h92;
		ram[15'h45A] = 8'h00;
		ram[15'h45B] = 8'h3E;
		ram[15'h45C] = 8'h07;
		ram[15'h45D] = 8'h21;
		ram[15'h45E] = 8'h06;
		ram[15'h45F] = 8'h05;
		ram[15'h460] = 8'hA7;
		ram[15'h461] = 8'hA7;
		ram[15'h462] = 8'hA7;
		ram[15'h463] = 8'hA0;
		ram[15'h464] = 8'hA7;
		ram[15'h465] = 8'hA1;
		ram[15'h466] = 8'hA7;
		ram[15'h467] = 8'hA2;
		ram[15'h468] = 8'hA7;
		ram[15'h469] = 8'hA3;
		ram[15'h46A] = 8'hA7;
		ram[15'h46B] = 8'hA4;
		ram[15'h46C] = 8'hA7;
		ram[15'h46D] = 8'hA5;
		ram[15'h46E] = 8'h21;
		ram[15'h46F] = 8'h92;
		ram[15'h470] = 8'h00;
		ram[15'h471] = 8'h36;
		ram[15'h472] = 8'h08;
		ram[15'h473] = 8'hA7;
		ram[15'h474] = 8'hA6;
		ram[15'h475] = 8'hA7;
		ram[15'h476] = 8'hDD;
		ram[15'h477] = 8'hA6;
		ram[15'h478] = 8'h00;
		ram[15'h479] = 8'hA7;
		ram[15'h47A] = 8'hFD;
		ram[15'h47B] = 8'hA6;
		ram[15'h47C] = 8'h01;
		ram[15'h47D] = 8'hA7;
		ram[15'h47E] = 8'hE6;
		ram[15'h47F] = 8'h0B;
		ram[15'h480] = 8'h32;
		ram[15'h481] = 8'h92;
		ram[15'h482] = 8'h00;
		ram[15'h483] = 8'h3E;
		ram[15'h484] = 8'h07;
		ram[15'h485] = 8'h21;
		ram[15'h486] = 8'h06;
		ram[15'h487] = 8'h05;
		ram[15'h488] = 8'hB7;
		ram[15'h489] = 8'hB7;
		ram[15'h48A] = 8'hB7;
		ram[15'h48B] = 8'hB0;
		ram[15'h48C] = 8'hB7;
		ram[15'h48D] = 8'hB1;
		ram[15'h48E] = 8'hB7;
		ram[15'h48F] = 8'hB2;
		ram[15'h490] = 8'hB7;
		ram[15'h491] = 8'hB3;
		ram[15'h492] = 8'hB7;
		ram[15'h493] = 8'hB4;
		ram[15'h494] = 8'hB7;
		ram[15'h495] = 8'hB5;
		ram[15'h496] = 8'h21;
		ram[15'h497] = 8'h92;
		ram[15'h498] = 8'h00;
		ram[15'h499] = 8'h36;
		ram[15'h49A] = 8'h08;
		ram[15'h49B] = 8'hB7;
		ram[15'h49C] = 8'hB6;
		ram[15'h49D] = 8'hB7;
		ram[15'h49E] = 8'hDD;
		ram[15'h49F] = 8'hB6;
		ram[15'h4A0] = 8'h00;
		ram[15'h4A1] = 8'hB7;
		ram[15'h4A2] = 8'hFD;
		ram[15'h4A3] = 8'hB6;
		ram[15'h4A4] = 8'h01;
		ram[15'h4A5] = 8'hB7;
		ram[15'h4A6] = 8'hF6;
		ram[15'h4A7] = 8'h0B;
		ram[15'h4A8] = 8'h32;
		ram[15'h4A9] = 8'h92;
		ram[15'h4AA] = 8'h00;
		ram[15'h4AB] = 8'h3E;
		ram[15'h4AC] = 8'h07;
		ram[15'h4AD] = 8'h21;
		ram[15'h4AE] = 8'h06;
		ram[15'h4AF] = 8'h05;
		ram[15'h4B0] = 8'hAF;
		ram[15'h4B1] = 8'hAF;
		ram[15'h4B2] = 8'hAF;
		ram[15'h4B3] = 8'hA8;
		ram[15'h4B4] = 8'hAF;
		ram[15'h4B5] = 8'hA9;
		ram[15'h4B6] = 8'hAF;
		ram[15'h4B7] = 8'hAA;
		ram[15'h4B8] = 8'hAF;
		ram[15'h4B9] = 8'hAB;
		ram[15'h4BA] = 8'hAF;
		ram[15'h4BB] = 8'hAC;
		ram[15'h4BC] = 8'hAF;
		ram[15'h4BD] = 8'hAD;
		ram[15'h4BE] = 8'h21;
		ram[15'h4BF] = 8'h92;
		ram[15'h4C0] = 8'h00;
		ram[15'h4C1] = 8'h36;
		ram[15'h4C2] = 8'h08;
		ram[15'h4C3] = 8'hAF;
		ram[15'h4C4] = 8'hAE;
		ram[15'h4C5] = 8'hAF;
		ram[15'h4C6] = 8'hDD;
		ram[15'h4C7] = 8'hAE;
		ram[15'h4C8] = 8'h00;
		ram[15'h4C9] = 8'hAF;
		ram[15'h4CA] = 8'hFD;
		ram[15'h4CB] = 8'hAE;
		ram[15'h4CC] = 8'h01;
		ram[15'h4CD] = 8'hAF;
		ram[15'h4CE] = 8'hEE;
		ram[15'h4CF] = 8'h0B;
		ram[15'h4D0] = 8'h32;
		ram[15'h4D1] = 8'h92;
		ram[15'h4D2] = 8'h00;
		ram[15'h4D3] = 8'h3E;
		ram[15'h4D4] = 8'h07;
		ram[15'h4D5] = 8'h21;
		ram[15'h4D6] = 8'h06;
		ram[15'h4D7] = 8'h05;
		ram[15'h4D8] = 8'hBF;
		ram[15'h4D9] = 8'hBF;
		ram[15'h4DA] = 8'hBF;
		ram[15'h4DB] = 8'hB8;
		ram[15'h4DC] = 8'hBF;
		ram[15'h4DD] = 8'hB9;
		ram[15'h4DE] = 8'hBF;
		ram[15'h4DF] = 8'hBA;
		ram[15'h4E0] = 8'hBF;
		ram[15'h4E1] = 8'hBB;
		ram[15'h4E2] = 8'hBF;
		ram[15'h4E3] = 8'hBC;
		ram[15'h4E4] = 8'hBF;
		ram[15'h4E5] = 8'hBD;
		ram[15'h4E6] = 8'h21;
		ram[15'h4E7] = 8'h92;
		ram[15'h4E8] = 8'h00;
		ram[15'h4E9] = 8'h36;
		ram[15'h4EA] = 8'h08;
		ram[15'h4EB] = 8'hBF;
		ram[15'h4EC] = 8'hBE;
		ram[15'h4ED] = 8'hBF;
		ram[15'h4EE] = 8'hDD;
		ram[15'h4EF] = 8'hBE;
		ram[15'h4F0] = 8'h00;
		ram[15'h4F1] = 8'hBF;
		ram[15'h4F2] = 8'hFD;
		ram[15'h4F3] = 8'hBE;
		ram[15'h4F4] = 8'h01;
		ram[15'h4F5] = 8'hBF;
		ram[15'h4F6] = 8'hFE;
		ram[15'h4F7] = 8'h0B;
		ram[15'h4F8] = 8'h32;
		ram[15'h4F9] = 8'h92;
		ram[15'h4FA] = 8'h00;
		ram[15'h4FB] = 8'hDD;
		ram[15'h4FC] = 8'h21;
		ram[15'h4FD] = 8'h92;
		ram[15'h4FE] = 8'h00;
		ram[15'h4FF] = 8'hFD;
		ram[15'h500] = 8'h21;
		ram[15'h501] = 8'h93;
		ram[15'h502] = 8'h00;
		ram[15'h503] = 8'h3E;
		ram[15'h504] = 8'h01;
		ram[15'h505] = 8'h3C;
		ram[15'h506] = 8'hDD;
		ram[15'h507] = 8'h77;
		ram[15'h508] = 8'h00;
		ram[15'h509] = 8'h47;
		ram[15'h50A] = 8'h04;
		ram[15'h50B] = 8'hDD;
		ram[15'h50C] = 8'h70;
		ram[15'h50D] = 8'h00;
		ram[15'h50E] = 8'h48;
		ram[15'h50F] = 8'h0C;
		ram[15'h510] = 8'hDD;
		ram[15'h511] = 8'h71;
		ram[15'h512] = 8'h00;
		ram[15'h513] = 8'h51;
		ram[15'h514] = 8'h14;
		ram[15'h515] = 8'hDD;
		ram[15'h516] = 8'h72;
		ram[15'h517] = 8'h00;
		ram[15'h518] = 8'h5A;
		ram[15'h519] = 8'h1C;
		ram[15'h51A] = 8'hDD;
		ram[15'h51B] = 8'h73;
		ram[15'h51C] = 8'h00;
		ram[15'h51D] = 8'h63;
		ram[15'h51E] = 8'h24;
		ram[15'h51F] = 8'hDD;
		ram[15'h520] = 8'h74;
		ram[15'h521] = 8'h00;
		ram[15'h522] = 8'h6C;
		ram[15'h523] = 8'h2C;
		ram[15'h524] = 8'hDD;
		ram[15'h525] = 8'h75;
		ram[15'h526] = 8'h00;
		ram[15'h527] = 8'hDD;
		ram[15'h528] = 8'h34;
		ram[15'h529] = 8'h00;
		ram[15'h52A] = 8'hDD;
		ram[15'h52B] = 8'h7E;
		ram[15'h52C] = 8'h00;
		ram[15'h52D] = 8'hFD;
		ram[15'h52E] = 8'h77;
		ram[15'h52F] = 8'h00;
		ram[15'h530] = 8'hFD;
		ram[15'h531] = 8'h34;
		ram[15'h532] = 8'h00;
		ram[15'h533] = 8'h21;
		ram[15'h534] = 8'h92;
		ram[15'h535] = 8'h00;
		ram[15'h536] = 8'h34;
		ram[15'h537] = 8'h3E;
		ram[15'h538] = 8'hFE;
		ram[15'h539] = 8'h3D;
		ram[15'h53A] = 8'hDD;
		ram[15'h53B] = 8'h77;
		ram[15'h53C] = 8'h00;
		ram[15'h53D] = 8'h47;
		ram[15'h53E] = 8'h05;
		ram[15'h53F] = 8'hDD;
		ram[15'h540] = 8'h70;
		ram[15'h541] = 8'h00;
		ram[15'h542] = 8'h48;
		ram[15'h543] = 8'h0D;
		ram[15'h544] = 8'hDD;
		ram[15'h545] = 8'h71;
		ram[15'h546] = 8'h00;
		ram[15'h547] = 8'h51;
		ram[15'h548] = 8'h15;
		ram[15'h549] = 8'hDD;
		ram[15'h54A] = 8'h72;
		ram[15'h54B] = 8'h00;
		ram[15'h54C] = 8'h5A;
		ram[15'h54D] = 8'h1D;
		ram[15'h54E] = 8'hDD;
		ram[15'h54F] = 8'h73;
		ram[15'h550] = 8'h00;
		ram[15'h551] = 8'h63;
		ram[15'h552] = 8'h25;
		ram[15'h553] = 8'hDD;
		ram[15'h554] = 8'h74;
		ram[15'h555] = 8'h00;
		ram[15'h556] = 8'h6C;
		ram[15'h557] = 8'h2D;
		ram[15'h558] = 8'hDD;
		ram[15'h559] = 8'h75;
		ram[15'h55A] = 8'h00;
		ram[15'h55B] = 8'hDD;
		ram[15'h55C] = 8'h35;
		ram[15'h55D] = 8'h00;
		ram[15'h55E] = 8'hDD;
		ram[15'h55F] = 8'h7E;
		ram[15'h560] = 8'h00;
		ram[15'h561] = 8'hFD;
		ram[15'h562] = 8'h77;
		ram[15'h563] = 8'h00;
		ram[15'h564] = 8'hFD;
		ram[15'h565] = 8'h35;
		ram[15'h566] = 8'h00;
		ram[15'h567] = 8'h21;
		ram[15'h568] = 8'h92;
		ram[15'h569] = 8'h00;
		ram[15'h56A] = 8'h35;
		ram[15'h56B] = 8'hC9;
		ram[15'h56C] = 8'h3E;
		ram[15'h56D] = 8'h0A;
		ram[15'h56E] = 8'hD3;
		ram[15'h56F] = 8'h01;
		ram[15'h570] = 8'h27;
		ram[15'h571] = 8'h2F;
		ram[15'h572] = 8'hED;
		ram[15'h573] = 8'h44;
		ram[15'h574] = 8'h3F;
		ram[15'h575] = 8'h37;
		ram[15'h576] = 8'h00;
		ram[15'h577] = 8'hF3;
		ram[15'h578] = 8'hED;
		ram[15'h579] = 8'h46;
		ram[15'h57A] = 8'hED;
		ram[15'h57B] = 8'h56;
		ram[15'h57C] = 8'hED;
		ram[15'h57D] = 8'h5E;
		ram[15'h57E] = 8'hED;
		ram[15'h57F] = 8'h46;
		ram[15'h580] = 8'hFB;
		ram[15'h581] = 8'hC9;
		ram[15'h582] = 8'h3E;
		ram[15'h583] = 8'h0B;
		ram[15'h584] = 8'hD3;
		ram[15'h585] = 8'h01;
		ram[15'h586] = 8'hC9;
		ram[15'h587] = 8'h3E;
		ram[15'h588] = 8'h0C;
		ram[15'h589] = 8'hD3;
		ram[15'h58A] = 8'h01;
		ram[15'h58B] = 8'h21;
		ram[15'h58C] = 8'h00;
		ram[15'h58D] = 8'h00;
		ram[15'h58E] = 8'h39;
		ram[15'h58F] = 8'h22;
		ram[15'h590] = 8'h96;
		ram[15'h591] = 8'h00;
		ram[15'h592] = 8'h21;
		ram[15'h593] = 8'h00;
		ram[15'h594] = 8'h00;
		ram[15'h595] = 8'h01;
		ram[15'h596] = 8'h01;
		ram[15'h597] = 8'h01;
		ram[15'h598] = 8'h09;
		ram[15'h599] = 8'h22;
		ram[15'h59A] = 8'h96;
		ram[15'h59B] = 8'h00;
		ram[15'h59C] = 8'h21;
		ram[15'h59D] = 8'h00;
		ram[15'h59E] = 8'h00;
		ram[15'h59F] = 8'h11;
		ram[15'h5A0] = 8'h02;
		ram[15'h5A1] = 8'h02;
		ram[15'h5A2] = 8'h19;
		ram[15'h5A3] = 8'h22;
		ram[15'h5A4] = 8'h96;
		ram[15'h5A5] = 8'h00;
		ram[15'h5A6] = 8'h21;
		ram[15'h5A7] = 8'h00;
		ram[15'h5A8] = 8'h00;
		ram[15'h5A9] = 8'h21;
		ram[15'h5AA] = 8'h03;
		ram[15'h5AB] = 8'h03;
		ram[15'h5AC] = 8'h29;
		ram[15'h5AD] = 8'h22;
		ram[15'h5AE] = 8'h96;
		ram[15'h5AF] = 8'h00;
		ram[15'h5B0] = 8'hDD;
		ram[15'h5B1] = 8'h21;
		ram[15'h5B2] = 8'h00;
		ram[15'h5B3] = 8'h00;
		ram[15'h5B4] = 8'hDD;
		ram[15'h5B5] = 8'h39;
		ram[15'h5B6] = 8'hDD;
		ram[15'h5B7] = 8'h22;
		ram[15'h5B8] = 8'h96;
		ram[15'h5B9] = 8'h00;
		ram[15'h5BA] = 8'hDD;
		ram[15'h5BB] = 8'h21;
		ram[15'h5BC] = 8'h00;
		ram[15'h5BD] = 8'h00;
		ram[15'h5BE] = 8'h01;
		ram[15'h5BF] = 8'h01;
		ram[15'h5C0] = 8'h01;
		ram[15'h5C1] = 8'hDD;
		ram[15'h5C2] = 8'h09;
		ram[15'h5C3] = 8'hDD;
		ram[15'h5C4] = 8'h22;
		ram[15'h5C5] = 8'h96;
		ram[15'h5C6] = 8'h00;
		ram[15'h5C7] = 8'hDD;
		ram[15'h5C8] = 8'h21;
		ram[15'h5C9] = 8'h00;
		ram[15'h5CA] = 8'h00;
		ram[15'h5CB] = 8'h11;
		ram[15'h5CC] = 8'h02;
		ram[15'h5CD] = 8'h02;
		ram[15'h5CE] = 8'hDD;
		ram[15'h5CF] = 8'h19;
		ram[15'h5D0] = 8'hDD;
		ram[15'h5D1] = 8'h22;
		ram[15'h5D2] = 8'h96;
		ram[15'h5D3] = 8'h00;
		ram[15'h5D4] = 8'hDD;
		ram[15'h5D5] = 8'h21;
		ram[15'h5D6] = 8'h00;
		ram[15'h5D7] = 8'h00;
		ram[15'h5D8] = 8'hDD;
		ram[15'h5D9] = 8'h21;
		ram[15'h5DA] = 8'h03;
		ram[15'h5DB] = 8'h03;
		ram[15'h5DC] = 8'hDD;
		ram[15'h5DD] = 8'h29;
		ram[15'h5DE] = 8'hDD;
		ram[15'h5DF] = 8'h22;
		ram[15'h5E0] = 8'h96;
		ram[15'h5E1] = 8'h00;
		ram[15'h5E2] = 8'hFD;
		ram[15'h5E3] = 8'h21;
		ram[15'h5E4] = 8'h00;
		ram[15'h5E5] = 8'h00;
		ram[15'h5E6] = 8'hFD;
		ram[15'h5E7] = 8'h39;
		ram[15'h5E8] = 8'hFD;
		ram[15'h5E9] = 8'h22;
		ram[15'h5EA] = 8'h96;
		ram[15'h5EB] = 8'h00;
		ram[15'h5EC] = 8'hFD;
		ram[15'h5ED] = 8'h21;
		ram[15'h5EE] = 8'h00;
		ram[15'h5EF] = 8'h00;
		ram[15'h5F0] = 8'h01;
		ram[15'h5F1] = 8'h01;
		ram[15'h5F2] = 8'h01;
		ram[15'h5F3] = 8'hFD;
		ram[15'h5F4] = 8'h09;
		ram[15'h5F5] = 8'hFD;
		ram[15'h5F6] = 8'h22;
		ram[15'h5F7] = 8'h96;
		ram[15'h5F8] = 8'h00;
		ram[15'h5F9] = 8'hFD;
		ram[15'h5FA] = 8'h21;
		ram[15'h5FB] = 8'h00;
		ram[15'h5FC] = 8'h00;
		ram[15'h5FD] = 8'h11;
		ram[15'h5FE] = 8'h02;
		ram[15'h5FF] = 8'h02;
		ram[15'h600] = 8'hFD;
		ram[15'h601] = 8'h19;
		ram[15'h602] = 8'hFD;
		ram[15'h603] = 8'h22;
		ram[15'h604] = 8'h96;
		ram[15'h605] = 8'h00;
		ram[15'h606] = 8'hFD;
		ram[15'h607] = 8'h21;
		ram[15'h608] = 8'h00;
		ram[15'h609] = 8'h00;
		ram[15'h60A] = 8'hFD;
		ram[15'h60B] = 8'h21;
		ram[15'h60C] = 8'h03;
		ram[15'h60D] = 8'h03;
		ram[15'h60E] = 8'hFD;
		ram[15'h60F] = 8'h29;
		ram[15'h610] = 8'hFD;
		ram[15'h611] = 8'h22;
		ram[15'h612] = 8'h96;
		ram[15'h613] = 8'h00;
		ram[15'h614] = 8'h21;
		ram[15'h615] = 8'h02;
		ram[15'h616] = 8'h01;
		ram[15'h617] = 8'h11;
		ram[15'h618] = 8'h04;
		ram[15'h619] = 8'h03;
		ram[15'h61A] = 8'h01;
		ram[15'h61B] = 8'h06;
		ram[15'h61C] = 8'h05;
		ram[15'h61D] = 8'hDD;
		ram[15'h61E] = 8'h21;
		ram[15'h61F] = 8'h08;
		ram[15'h620] = 8'h07;
		ram[15'h621] = 8'hFD;
		ram[15'h622] = 8'h21;
		ram[15'h623] = 8'h0A;
		ram[15'h624] = 8'h09;
		ram[15'h625] = 8'h23;
		ram[15'h626] = 8'h22;
		ram[15'h627] = 8'h96;
		ram[15'h628] = 8'h00;
		ram[15'h629] = 8'hDD;
		ram[15'h62A] = 8'h23;
		ram[15'h62B] = 8'hDD;
		ram[15'h62C] = 8'h22;
		ram[15'h62D] = 8'h96;
		ram[15'h62E] = 8'h00;
		ram[15'h62F] = 8'hFD;
		ram[15'h630] = 8'h23;
		ram[15'h631] = 8'hFD;
		ram[15'h632] = 8'h22;
		ram[15'h633] = 8'h96;
		ram[15'h634] = 8'h00;
		ram[15'h635] = 8'h13;
		ram[15'h636] = 8'hED;
		ram[15'h637] = 8'h53;
		ram[15'h638] = 8'h96;
		ram[15'h639] = 8'h00;
		ram[15'h63A] = 8'h03;
		ram[15'h63B] = 8'hED;
		ram[15'h63C] = 8'h43;
		ram[15'h63D] = 8'h96;
		ram[15'h63E] = 8'h00;
		ram[15'h63F] = 8'h2B;
		ram[15'h640] = 8'h22;
		ram[15'h641] = 8'h96;
		ram[15'h642] = 8'h00;
		ram[15'h643] = 8'hDD;
		ram[15'h644] = 8'h2B;
		ram[15'h645] = 8'hDD;
		ram[15'h646] = 8'h22;
		ram[15'h647] = 8'h96;
		ram[15'h648] = 8'h00;
		ram[15'h649] = 8'hFD;
		ram[15'h64A] = 8'h2B;
		ram[15'h64B] = 8'hFD;
		ram[15'h64C] = 8'h22;
		ram[15'h64D] = 8'h96;
		ram[15'h64E] = 8'h00;
		ram[15'h64F] = 8'h1B;
		ram[15'h650] = 8'hED;
		ram[15'h651] = 8'h53;
		ram[15'h652] = 8'h96;
		ram[15'h653] = 8'h00;
		ram[15'h654] = 8'h0B;
		ram[15'h655] = 8'hED;
		ram[15'h656] = 8'h43;
		ram[15'h657] = 8'h96;
		ram[15'h658] = 8'h00;
		ram[15'h659] = 8'hC9;
		ram[15'h65A] = 8'h3E;
		ram[15'h65B] = 8'h0D;
		ram[15'h65C] = 8'hD3;
		ram[15'h65D] = 8'h01;
		ram[15'h65E] = 8'h3E;
		ram[15'h65F] = 8'hAA;
		ram[15'h660] = 8'h07;
		ram[15'h661] = 8'h17;
		ram[15'h662] = 8'h0F;
		ram[15'h663] = 8'h1F;
		ram[15'h664] = 8'hF5;
		ram[15'h665] = 8'hE5;
		ram[15'h666] = 8'hE1;
		ram[15'h667] = 8'hF1;
		ram[15'h668] = 8'h21;
		ram[15'h669] = 8'h96;
		ram[15'h66A] = 8'h00;
		ram[15'h66B] = 8'h36;
		ram[15'h66C] = 8'h08;
		ram[15'h66D] = 8'hE5;
		ram[15'h66E] = 8'hDD;
		ram[15'h66F] = 8'hE1;
		ram[15'h670] = 8'hDD;
		ram[15'h671] = 8'h36;
		ram[15'h672] = 8'h01;
		ram[15'h673] = 8'h09;
		ram[15'h674] = 8'hE5;
		ram[15'h675] = 8'hFD;
		ram[15'h676] = 8'hE1;
		ram[15'h677] = 8'hFD;
		ram[15'h678] = 8'h36;
		ram[15'h679] = 8'h02;
		ram[15'h67A] = 8'h0A;
		ram[15'h67B] = 8'h01;
		ram[15'h67C] = 8'h02;
		ram[15'h67D] = 8'h01;
		ram[15'h67E] = 8'h11;
		ram[15'h67F] = 8'h04;
		ram[15'h680] = 8'h03;
		ram[15'h681] = 8'h21;
		ram[15'h682] = 8'h06;
		ram[15'h683] = 8'h05;
		ram[15'h684] = 8'h3E;
		ram[15'h685] = 8'h07;
		ram[15'h686] = 8'h21;
		ram[15'h687] = 8'h06;
		ram[15'h688] = 8'h05;
		ram[15'h689] = 8'hCB;
		ram[15'h68A] = 8'h00;
		ram[15'h68B] = 8'hCB;
		ram[15'h68C] = 8'h01;
		ram[15'h68D] = 8'hCB;
		ram[15'h68E] = 8'h02;
		ram[15'h68F] = 8'hCB;
		ram[15'h690] = 8'h03;
		ram[15'h691] = 8'hCB;
		ram[15'h692] = 8'h04;
		ram[15'h693] = 8'hCB;
		ram[15'h694] = 8'h05;
		ram[15'h695] = 8'hCB;
		ram[15'h696] = 8'h07;
		ram[15'h697] = 8'h21;
		ram[15'h698] = 8'h96;
		ram[15'h699] = 8'h00;
		ram[15'h69A] = 8'hCB;
		ram[15'h69B] = 8'h06;
		ram[15'h69C] = 8'hDD;
		ram[15'h69D] = 8'hCB;
		ram[15'h69E] = 8'h01;
		ram[15'h69F] = 8'h06;
		ram[15'h6A0] = 8'hDD;
		ram[15'h6A1] = 8'hCB;
		ram[15'h6A2] = 8'h02;
		ram[15'h6A3] = 8'h06;
		ram[15'h6A4] = 8'h21;
		ram[15'h6A5] = 8'h06;
		ram[15'h6A6] = 8'h05;
		ram[15'h6A7] = 8'hCB;
		ram[15'h6A8] = 8'h08;
		ram[15'h6A9] = 8'hCB;
		ram[15'h6AA] = 8'h09;
		ram[15'h6AB] = 8'hCB;
		ram[15'h6AC] = 8'h0A;
		ram[15'h6AD] = 8'hCB;
		ram[15'h6AE] = 8'h0B;
		ram[15'h6AF] = 8'hCB;
		ram[15'h6B0] = 8'h0C;
		ram[15'h6B1] = 8'hCB;
		ram[15'h6B2] = 8'h0D;
		ram[15'h6B3] = 8'hCB;
		ram[15'h6B4] = 8'h0F;
		ram[15'h6B5] = 8'h21;
		ram[15'h6B6] = 8'h96;
		ram[15'h6B7] = 8'h00;
		ram[15'h6B8] = 8'hCB;
		ram[15'h6B9] = 8'h0E;
		ram[15'h6BA] = 8'hDD;
		ram[15'h6BB] = 8'hCB;
		ram[15'h6BC] = 8'h01;
		ram[15'h6BD] = 8'h0E;
		ram[15'h6BE] = 8'hDD;
		ram[15'h6BF] = 8'hCB;
		ram[15'h6C0] = 8'h02;
		ram[15'h6C1] = 8'h0E;
		ram[15'h6C2] = 8'h21;
		ram[15'h6C3] = 8'h06;
		ram[15'h6C4] = 8'h05;
		ram[15'h6C5] = 8'hCB;
		ram[15'h6C6] = 8'h10;
		ram[15'h6C7] = 8'hCB;
		ram[15'h6C8] = 8'h11;
		ram[15'h6C9] = 8'hCB;
		ram[15'h6CA] = 8'h12;
		ram[15'h6CB] = 8'hCB;
		ram[15'h6CC] = 8'h13;
		ram[15'h6CD] = 8'hCB;
		ram[15'h6CE] = 8'h14;
		ram[15'h6CF] = 8'hCB;
		ram[15'h6D0] = 8'h15;
		ram[15'h6D1] = 8'hCB;
		ram[15'h6D2] = 8'h17;
		ram[15'h6D3] = 8'h21;
		ram[15'h6D4] = 8'h96;
		ram[15'h6D5] = 8'h00;
		ram[15'h6D6] = 8'hCB;
		ram[15'h6D7] = 8'h16;
		ram[15'h6D8] = 8'hDD;
		ram[15'h6D9] = 8'hCB;
		ram[15'h6DA] = 8'h01;
		ram[15'h6DB] = 8'h16;
		ram[15'h6DC] = 8'hDD;
		ram[15'h6DD] = 8'hCB;
		ram[15'h6DE] = 8'h02;
		ram[15'h6DF] = 8'h16;
		ram[15'h6E0] = 8'h21;
		ram[15'h6E1] = 8'h06;
		ram[15'h6E2] = 8'h05;
		ram[15'h6E3] = 8'hCB;
		ram[15'h6E4] = 8'h18;
		ram[15'h6E5] = 8'hCB;
		ram[15'h6E6] = 8'h19;
		ram[15'h6E7] = 8'hCB;
		ram[15'h6E8] = 8'h1A;
		ram[15'h6E9] = 8'hCB;
		ram[15'h6EA] = 8'h1B;
		ram[15'h6EB] = 8'hCB;
		ram[15'h6EC] = 8'h1C;
		ram[15'h6ED] = 8'hCB;
		ram[15'h6EE] = 8'h1D;
		ram[15'h6EF] = 8'hCB;
		ram[15'h6F0] = 8'h1F;
		ram[15'h6F1] = 8'h21;
		ram[15'h6F2] = 8'h96;
		ram[15'h6F3] = 8'h00;
		ram[15'h6F4] = 8'hCB;
		ram[15'h6F5] = 8'h1E;
		ram[15'h6F6] = 8'hDD;
		ram[15'h6F7] = 8'hCB;
		ram[15'h6F8] = 8'h01;
		ram[15'h6F9] = 8'h1E;
		ram[15'h6FA] = 8'hDD;
		ram[15'h6FB] = 8'hCB;
		ram[15'h6FC] = 8'h02;
		ram[15'h6FD] = 8'h1E;
		ram[15'h6FE] = 8'h21;
		ram[15'h6FF] = 8'h06;
		ram[15'h700] = 8'h05;
		ram[15'h701] = 8'hCB;
		ram[15'h702] = 8'h20;
		ram[15'h703] = 8'hCB;
		ram[15'h704] = 8'h21;
		ram[15'h705] = 8'hCB;
		ram[15'h706] = 8'h22;
		ram[15'h707] = 8'hCB;
		ram[15'h708] = 8'h23;
		ram[15'h709] = 8'hCB;
		ram[15'h70A] = 8'h24;
		ram[15'h70B] = 8'hCB;
		ram[15'h70C] = 8'h25;
		ram[15'h70D] = 8'hCB;
		ram[15'h70E] = 8'h27;
		ram[15'h70F] = 8'h21;
		ram[15'h710] = 8'h96;
		ram[15'h711] = 8'h00;
		ram[15'h712] = 8'hCB;
		ram[15'h713] = 8'h26;
		ram[15'h714] = 8'hDD;
		ram[15'h715] = 8'hCB;
		ram[15'h716] = 8'h01;
		ram[15'h717] = 8'h26;
		ram[15'h718] = 8'hDD;
		ram[15'h719] = 8'hCB;
		ram[15'h71A] = 8'h02;
		ram[15'h71B] = 8'h26;
		ram[15'h71C] = 8'h21;
		ram[15'h71D] = 8'h06;
		ram[15'h71E] = 8'h05;
		ram[15'h71F] = 8'hCB;
		ram[15'h720] = 8'h28;
		ram[15'h721] = 8'hCB;
		ram[15'h722] = 8'h29;
		ram[15'h723] = 8'hCB;
		ram[15'h724] = 8'h2A;
		ram[15'h725] = 8'hCB;
		ram[15'h726] = 8'h2B;
		ram[15'h727] = 8'hCB;
		ram[15'h728] = 8'h2C;
		ram[15'h729] = 8'hCB;
		ram[15'h72A] = 8'h2D;
		ram[15'h72B] = 8'hCB;
		ram[15'h72C] = 8'h2F;
		ram[15'h72D] = 8'h21;
		ram[15'h72E] = 8'h96;
		ram[15'h72F] = 8'h00;
		ram[15'h730] = 8'hCB;
		ram[15'h731] = 8'h2E;
		ram[15'h732] = 8'hDD;
		ram[15'h733] = 8'hCB;
		ram[15'h734] = 8'h01;
		ram[15'h735] = 8'h2E;
		ram[15'h736] = 8'hDD;
		ram[15'h737] = 8'hCB;
		ram[15'h738] = 8'h02;
		ram[15'h739] = 8'h2E;
		ram[15'h73A] = 8'h21;
		ram[15'h73B] = 8'h06;
		ram[15'h73C] = 8'h05;
		ram[15'h73D] = 8'hCB;
		ram[15'h73E] = 8'h30;
		ram[15'h73F] = 8'hCB;
		ram[15'h740] = 8'h31;
		ram[15'h741] = 8'hCB;
		ram[15'h742] = 8'h32;
		ram[15'h743] = 8'hCB;
		ram[15'h744] = 8'h33;
		ram[15'h745] = 8'hCB;
		ram[15'h746] = 8'h34;
		ram[15'h747] = 8'hCB;
		ram[15'h748] = 8'h35;
		ram[15'h749] = 8'hCB;
		ram[15'h74A] = 8'h37;
		ram[15'h74B] = 8'h21;
		ram[15'h74C] = 8'h96;
		ram[15'h74D] = 8'h00;
		ram[15'h74E] = 8'hCB;
		ram[15'h74F] = 8'h36;
		ram[15'h750] = 8'hDD;
		ram[15'h751] = 8'hCB;
		ram[15'h752] = 8'h01;
		ram[15'h753] = 8'h36;
		ram[15'h754] = 8'hDD;
		ram[15'h755] = 8'hCB;
		ram[15'h756] = 8'h02;
		ram[15'h757] = 8'h36;
		ram[15'h758] = 8'h21;
		ram[15'h759] = 8'h06;
		ram[15'h75A] = 8'h05;
		ram[15'h75B] = 8'hCB;
		ram[15'h75C] = 8'h38;
		ram[15'h75D] = 8'hCB;
		ram[15'h75E] = 8'h39;
		ram[15'h75F] = 8'hCB;
		ram[15'h760] = 8'h3A;
		ram[15'h761] = 8'hCB;
		ram[15'h762] = 8'h3B;
		ram[15'h763] = 8'hCB;
		ram[15'h764] = 8'h3C;
		ram[15'h765] = 8'hCB;
		ram[15'h766] = 8'h3D;
		ram[15'h767] = 8'hCB;
		ram[15'h768] = 8'h3F;
		ram[15'h769] = 8'h21;
		ram[15'h76A] = 8'h96;
		ram[15'h76B] = 8'h00;
		ram[15'h76C] = 8'hCB;
		ram[15'h76D] = 8'h3E;
		ram[15'h76E] = 8'hDD;
		ram[15'h76F] = 8'hCB;
		ram[15'h770] = 8'h01;
		ram[15'h771] = 8'h3E;
		ram[15'h772] = 8'hDD;
		ram[15'h773] = 8'hCB;
		ram[15'h774] = 8'h02;
		ram[15'h775] = 8'h3E;
		ram[15'h776] = 8'hED;
		ram[15'h777] = 8'h6F;
		ram[15'h778] = 8'hED;
		ram[15'h779] = 8'h67;
		ram[15'h77A] = 8'hC9;
		ram[15'h77B] = 8'h3E;
		ram[15'h77C] = 8'h0E;
		ram[15'h77D] = 8'hD3;
		ram[15'h77E] = 8'h01;
		ram[15'h77F] = 8'h21;
		ram[15'h780] = 8'h96;
		ram[15'h781] = 8'h00;
		ram[15'h782] = 8'h36;
		ram[15'h783] = 8'h08;
		ram[15'h784] = 8'hE5;
		ram[15'h785] = 8'hDD;
		ram[15'h786] = 8'hE1;
		ram[15'h787] = 8'hDD;
		ram[15'h788] = 8'h36;
		ram[15'h789] = 8'h01;
		ram[15'h78A] = 8'h09;
		ram[15'h78B] = 8'hE5;
		ram[15'h78C] = 8'hFD;
		ram[15'h78D] = 8'hE1;
		ram[15'h78E] = 8'hFD;
		ram[15'h78F] = 8'h36;
		ram[15'h790] = 8'h02;
		ram[15'h791] = 8'h0A;
		ram[15'h792] = 8'h01;
		ram[15'h793] = 8'h02;
		ram[15'h794] = 8'h01;
		ram[15'h795] = 8'h11;
		ram[15'h796] = 8'h04;
		ram[15'h797] = 8'h03;
		ram[15'h798] = 8'h21;
		ram[15'h799] = 8'h06;
		ram[15'h79A] = 8'h05;
		ram[15'h79B] = 8'h3E;
		ram[15'h79C] = 8'h07;
		ram[15'h79D] = 8'h21;
		ram[15'h79E] = 8'h06;
		ram[15'h79F] = 8'h05;
		ram[15'h7A0] = 8'hCB;
		ram[15'h7A1] = 8'h40;
		ram[15'h7A2] = 8'hCB;
		ram[15'h7A3] = 8'h41;
		ram[15'h7A4] = 8'hCB;
		ram[15'h7A5] = 8'h42;
		ram[15'h7A6] = 8'hCB;
		ram[15'h7A7] = 8'h43;
		ram[15'h7A8] = 8'hCB;
		ram[15'h7A9] = 8'h44;
		ram[15'h7AA] = 8'hCB;
		ram[15'h7AB] = 8'h45;
		ram[15'h7AC] = 8'hCB;
		ram[15'h7AD] = 8'h47;
		ram[15'h7AE] = 8'h21;
		ram[15'h7AF] = 8'h96;
		ram[15'h7B0] = 8'h00;
		ram[15'h7B1] = 8'hCB;
		ram[15'h7B2] = 8'h46;
		ram[15'h7B3] = 8'hDD;
		ram[15'h7B4] = 8'hCB;
		ram[15'h7B5] = 8'h01;
		ram[15'h7B6] = 8'h46;
		ram[15'h7B7] = 8'hFD;
		ram[15'h7B8] = 8'hCB;
		ram[15'h7B9] = 8'h02;
		ram[15'h7BA] = 8'h46;
		ram[15'h7BB] = 8'h21;
		ram[15'h7BC] = 8'h06;
		ram[15'h7BD] = 8'h05;
		ram[15'h7BE] = 8'hCB;
		ram[15'h7BF] = 8'hC0;
		ram[15'h7C0] = 8'hCB;
		ram[15'h7C1] = 8'hC1;
		ram[15'h7C2] = 8'hCB;
		ram[15'h7C3] = 8'hC2;
		ram[15'h7C4] = 8'hCB;
		ram[15'h7C5] = 8'hC3;
		ram[15'h7C6] = 8'hCB;
		ram[15'h7C7] = 8'hC4;
		ram[15'h7C8] = 8'hCB;
		ram[15'h7C9] = 8'hC5;
		ram[15'h7CA] = 8'hCB;
		ram[15'h7CB] = 8'hC7;
		ram[15'h7CC] = 8'h21;
		ram[15'h7CD] = 8'h96;
		ram[15'h7CE] = 8'h00;
		ram[15'h7CF] = 8'hCB;
		ram[15'h7D0] = 8'hC6;
		ram[15'h7D1] = 8'hDD;
		ram[15'h7D2] = 8'hCB;
		ram[15'h7D3] = 8'h01;
		ram[15'h7D4] = 8'hC6;
		ram[15'h7D5] = 8'hFD;
		ram[15'h7D6] = 8'hCB;
		ram[15'h7D7] = 8'h02;
		ram[15'h7D8] = 8'hC6;
		ram[15'h7D9] = 8'h21;
		ram[15'h7DA] = 8'h06;
		ram[15'h7DB] = 8'h05;
		ram[15'h7DC] = 8'hCB;
		ram[15'h7DD] = 8'h80;
		ram[15'h7DE] = 8'hCB;
		ram[15'h7DF] = 8'h81;
		ram[15'h7E0] = 8'hCB;
		ram[15'h7E1] = 8'h82;
		ram[15'h7E2] = 8'hCB;
		ram[15'h7E3] = 8'h83;
		ram[15'h7E4] = 8'hCB;
		ram[15'h7E5] = 8'h84;
		ram[15'h7E6] = 8'hCB;
		ram[15'h7E7] = 8'h85;
		ram[15'h7E8] = 8'hCB;
		ram[15'h7E9] = 8'h87;
		ram[15'h7EA] = 8'h21;
		ram[15'h7EB] = 8'h96;
		ram[15'h7EC] = 8'h00;
		ram[15'h7ED] = 8'hCB;
		ram[15'h7EE] = 8'h86;
		ram[15'h7EF] = 8'hDD;
		ram[15'h7F0] = 8'hCB;
		ram[15'h7F1] = 8'h01;
		ram[15'h7F2] = 8'h86;
		ram[15'h7F3] = 8'hFD;
		ram[15'h7F4] = 8'hCB;
		ram[15'h7F5] = 8'h02;
		ram[15'h7F6] = 8'h86;
		ram[15'h7F7] = 8'h21;
		ram[15'h7F8] = 8'h06;
		ram[15'h7F9] = 8'h05;
		ram[15'h7FA] = 8'hCB;
		ram[15'h7FB] = 8'h48;
		ram[15'h7FC] = 8'hCB;
		ram[15'h7FD] = 8'h49;
		ram[15'h7FE] = 8'hCB;
		ram[15'h7FF] = 8'h4A;
		ram[15'h800] = 8'hCB;
		ram[15'h801] = 8'h4B;
		ram[15'h802] = 8'hCB;
		ram[15'h803] = 8'h4C;
		ram[15'h804] = 8'hCB;
		ram[15'h805] = 8'h4D;
		ram[15'h806] = 8'hCB;
		ram[15'h807] = 8'h4F;
		ram[15'h808] = 8'h21;
		ram[15'h809] = 8'h96;
		ram[15'h80A] = 8'h00;
		ram[15'h80B] = 8'hCB;
		ram[15'h80C] = 8'h4E;
		ram[15'h80D] = 8'hDD;
		ram[15'h80E] = 8'hCB;
		ram[15'h80F] = 8'h01;
		ram[15'h810] = 8'h4E;
		ram[15'h811] = 8'hFD;
		ram[15'h812] = 8'hCB;
		ram[15'h813] = 8'h02;
		ram[15'h814] = 8'h4E;
		ram[15'h815] = 8'h21;
		ram[15'h816] = 8'h06;
		ram[15'h817] = 8'h05;
		ram[15'h818] = 8'hCB;
		ram[15'h819] = 8'hC8;
		ram[15'h81A] = 8'hCB;
		ram[15'h81B] = 8'hC9;
		ram[15'h81C] = 8'hCB;
		ram[15'h81D] = 8'hCA;
		ram[15'h81E] = 8'hCB;
		ram[15'h81F] = 8'hCB;
		ram[15'h820] = 8'hCB;
		ram[15'h821] = 8'hCC;
		ram[15'h822] = 8'hCB;
		ram[15'h823] = 8'hCD;
		ram[15'h824] = 8'hCB;
		ram[15'h825] = 8'hCF;
		ram[15'h826] = 8'h21;
		ram[15'h827] = 8'h96;
		ram[15'h828] = 8'h00;
		ram[15'h829] = 8'hCB;
		ram[15'h82A] = 8'hCE;
		ram[15'h82B] = 8'hDD;
		ram[15'h82C] = 8'hCB;
		ram[15'h82D] = 8'h01;
		ram[15'h82E] = 8'hCE;
		ram[15'h82F] = 8'hFD;
		ram[15'h830] = 8'hCB;
		ram[15'h831] = 8'h02;
		ram[15'h832] = 8'hCE;
		ram[15'h833] = 8'h21;
		ram[15'h834] = 8'h06;
		ram[15'h835] = 8'h05;
		ram[15'h836] = 8'hCB;
		ram[15'h837] = 8'h88;
		ram[15'h838] = 8'hCB;
		ram[15'h839] = 8'h89;
		ram[15'h83A] = 8'hCB;
		ram[15'h83B] = 8'h8A;
		ram[15'h83C] = 8'hCB;
		ram[15'h83D] = 8'h8B;
		ram[15'h83E] = 8'hCB;
		ram[15'h83F] = 8'h8C;
		ram[15'h840] = 8'hCB;
		ram[15'h841] = 8'h8D;
		ram[15'h842] = 8'hCB;
		ram[15'h843] = 8'h8F;
		ram[15'h844] = 8'h21;
		ram[15'h845] = 8'h96;
		ram[15'h846] = 8'h00;
		ram[15'h847] = 8'hCB;
		ram[15'h848] = 8'h8E;
		ram[15'h849] = 8'hDD;
		ram[15'h84A] = 8'hCB;
		ram[15'h84B] = 8'h01;
		ram[15'h84C] = 8'h8E;
		ram[15'h84D] = 8'hFD;
		ram[15'h84E] = 8'hCB;
		ram[15'h84F] = 8'h02;
		ram[15'h850] = 8'h8E;
		ram[15'h851] = 8'h21;
		ram[15'h852] = 8'h06;
		ram[15'h853] = 8'h05;
		ram[15'h854] = 8'hCB;
		ram[15'h855] = 8'h50;
		ram[15'h856] = 8'hCB;
		ram[15'h857] = 8'h51;
		ram[15'h858] = 8'hCB;
		ram[15'h859] = 8'h52;
		ram[15'h85A] = 8'hCB;
		ram[15'h85B] = 8'h53;
		ram[15'h85C] = 8'hCB;
		ram[15'h85D] = 8'h54;
		ram[15'h85E] = 8'hCB;
		ram[15'h85F] = 8'h55;
		ram[15'h860] = 8'hCB;
		ram[15'h861] = 8'h57;
		ram[15'h862] = 8'h21;
		ram[15'h863] = 8'h96;
		ram[15'h864] = 8'h00;
		ram[15'h865] = 8'hCB;
		ram[15'h866] = 8'h56;
		ram[15'h867] = 8'hDD;
		ram[15'h868] = 8'hCB;
		ram[15'h869] = 8'h01;
		ram[15'h86A] = 8'h56;
		ram[15'h86B] = 8'hFD;
		ram[15'h86C] = 8'hCB;
		ram[15'h86D] = 8'h02;
		ram[15'h86E] = 8'h56;
		ram[15'h86F] = 8'h21;
		ram[15'h870] = 8'h06;
		ram[15'h871] = 8'h05;
		ram[15'h872] = 8'hCB;
		ram[15'h873] = 8'hD0;
		ram[15'h874] = 8'hCB;
		ram[15'h875] = 8'hD1;
		ram[15'h876] = 8'hCB;
		ram[15'h877] = 8'hD2;
		ram[15'h878] = 8'hCB;
		ram[15'h879] = 8'hD3;
		ram[15'h87A] = 8'hCB;
		ram[15'h87B] = 8'hD4;
		ram[15'h87C] = 8'hCB;
		ram[15'h87D] = 8'hD5;
		ram[15'h87E] = 8'hCB;
		ram[15'h87F] = 8'hD7;
		ram[15'h880] = 8'h21;
		ram[15'h881] = 8'h96;
		ram[15'h882] = 8'h00;
		ram[15'h883] = 8'hCB;
		ram[15'h884] = 8'hD6;
		ram[15'h885] = 8'hDD;
		ram[15'h886] = 8'hCB;
		ram[15'h887] = 8'h01;
		ram[15'h888] = 8'hD6;
		ram[15'h889] = 8'hFD;
		ram[15'h88A] = 8'hCB;
		ram[15'h88B] = 8'h02;
		ram[15'h88C] = 8'hD6;
		ram[15'h88D] = 8'h21;
		ram[15'h88E] = 8'h06;
		ram[15'h88F] = 8'h05;
		ram[15'h890] = 8'hCB;
		ram[15'h891] = 8'h90;
		ram[15'h892] = 8'hCB;
		ram[15'h893] = 8'h91;
		ram[15'h894] = 8'hCB;
		ram[15'h895] = 8'h92;
		ram[15'h896] = 8'hCB;
		ram[15'h897] = 8'h93;
		ram[15'h898] = 8'hCB;
		ram[15'h899] = 8'h94;
		ram[15'h89A] = 8'hCB;
		ram[15'h89B] = 8'h95;
		ram[15'h89C] = 8'hCB;
		ram[15'h89D] = 8'h97;
		ram[15'h89E] = 8'h21;
		ram[15'h89F] = 8'h96;
		ram[15'h8A0] = 8'h00;
		ram[15'h8A1] = 8'hCB;
		ram[15'h8A2] = 8'h96;
		ram[15'h8A3] = 8'hDD;
		ram[15'h8A4] = 8'hCB;
		ram[15'h8A5] = 8'h01;
		ram[15'h8A6] = 8'h96;
		ram[15'h8A7] = 8'hFD;
		ram[15'h8A8] = 8'hCB;
		ram[15'h8A9] = 8'h02;
		ram[15'h8AA] = 8'h96;
		ram[15'h8AB] = 8'h21;
		ram[15'h8AC] = 8'h06;
		ram[15'h8AD] = 8'h05;
		ram[15'h8AE] = 8'hCB;
		ram[15'h8AF] = 8'h58;
		ram[15'h8B0] = 8'hCB;
		ram[15'h8B1] = 8'h59;
		ram[15'h8B2] = 8'hCB;
		ram[15'h8B3] = 8'h5A;
		ram[15'h8B4] = 8'hCB;
		ram[15'h8B5] = 8'h5B;
		ram[15'h8B6] = 8'hCB;
		ram[15'h8B7] = 8'h5C;
		ram[15'h8B8] = 8'hCB;
		ram[15'h8B9] = 8'h5D;
		ram[15'h8BA] = 8'hCB;
		ram[15'h8BB] = 8'h5F;
		ram[15'h8BC] = 8'h21;
		ram[15'h8BD] = 8'h96;
		ram[15'h8BE] = 8'h00;
		ram[15'h8BF] = 8'hCB;
		ram[15'h8C0] = 8'h5E;
		ram[15'h8C1] = 8'hDD;
		ram[15'h8C2] = 8'hCB;
		ram[15'h8C3] = 8'h01;
		ram[15'h8C4] = 8'h5E;
		ram[15'h8C5] = 8'hFD;
		ram[15'h8C6] = 8'hCB;
		ram[15'h8C7] = 8'h02;
		ram[15'h8C8] = 8'h5E;
		ram[15'h8C9] = 8'h21;
		ram[15'h8CA] = 8'h06;
		ram[15'h8CB] = 8'h05;
		ram[15'h8CC] = 8'hCB;
		ram[15'h8CD] = 8'hD8;
		ram[15'h8CE] = 8'hCB;
		ram[15'h8CF] = 8'hD9;
		ram[15'h8D0] = 8'hCB;
		ram[15'h8D1] = 8'hDA;
		ram[15'h8D2] = 8'hCB;
		ram[15'h8D3] = 8'hDB;
		ram[15'h8D4] = 8'hCB;
		ram[15'h8D5] = 8'hDC;
		ram[15'h8D6] = 8'hCB;
		ram[15'h8D7] = 8'hDD;
		ram[15'h8D8] = 8'hCB;
		ram[15'h8D9] = 8'hDF;
		ram[15'h8DA] = 8'h21;
		ram[15'h8DB] = 8'h96;
		ram[15'h8DC] = 8'h00;
		ram[15'h8DD] = 8'hCB;
		ram[15'h8DE] = 8'hDE;
		ram[15'h8DF] = 8'hDD;
		ram[15'h8E0] = 8'hCB;
		ram[15'h8E1] = 8'h01;
		ram[15'h8E2] = 8'hDE;
		ram[15'h8E3] = 8'hFD;
		ram[15'h8E4] = 8'hCB;
		ram[15'h8E5] = 8'h02;
		ram[15'h8E6] = 8'hDE;
		ram[15'h8E7] = 8'h21;
		ram[15'h8E8] = 8'h06;
		ram[15'h8E9] = 8'h05;
		ram[15'h8EA] = 8'hCB;
		ram[15'h8EB] = 8'h98;
		ram[15'h8EC] = 8'hCB;
		ram[15'h8ED] = 8'h99;
		ram[15'h8EE] = 8'hCB;
		ram[15'h8EF] = 8'h9A;
		ram[15'h8F0] = 8'hCB;
		ram[15'h8F1] = 8'h9B;
		ram[15'h8F2] = 8'hCB;
		ram[15'h8F3] = 8'h9C;
		ram[15'h8F4] = 8'hCB;
		ram[15'h8F5] = 8'h9D;
		ram[15'h8F6] = 8'hCB;
		ram[15'h8F7] = 8'h9F;
		ram[15'h8F8] = 8'h21;
		ram[15'h8F9] = 8'h96;
		ram[15'h8FA] = 8'h00;
		ram[15'h8FB] = 8'hCB;
		ram[15'h8FC] = 8'h9E;
		ram[15'h8FD] = 8'hDD;
		ram[15'h8FE] = 8'hCB;
		ram[15'h8FF] = 8'h01;
		ram[15'h900] = 8'h9E;
		ram[15'h901] = 8'hFD;
		ram[15'h902] = 8'hCB;
		ram[15'h903] = 8'h02;
		ram[15'h904] = 8'h9E;
		ram[15'h905] = 8'h21;
		ram[15'h906] = 8'h06;
		ram[15'h907] = 8'h05;
		ram[15'h908] = 8'hCB;
		ram[15'h909] = 8'h60;
		ram[15'h90A] = 8'hCB;
		ram[15'h90B] = 8'h61;
		ram[15'h90C] = 8'hCB;
		ram[15'h90D] = 8'h62;
		ram[15'h90E] = 8'hCB;
		ram[15'h90F] = 8'h63;
		ram[15'h910] = 8'hCB;
		ram[15'h911] = 8'h64;
		ram[15'h912] = 8'hCB;
		ram[15'h913] = 8'h65;
		ram[15'h914] = 8'hCB;
		ram[15'h915] = 8'h67;
		ram[15'h916] = 8'h21;
		ram[15'h917] = 8'h96;
		ram[15'h918] = 8'h00;
		ram[15'h919] = 8'hCB;
		ram[15'h91A] = 8'h66;
		ram[15'h91B] = 8'hDD;
		ram[15'h91C] = 8'hCB;
		ram[15'h91D] = 8'h01;
		ram[15'h91E] = 8'h66;
		ram[15'h91F] = 8'hFD;
		ram[15'h920] = 8'hCB;
		ram[15'h921] = 8'h02;
		ram[15'h922] = 8'h66;
		ram[15'h923] = 8'h21;
		ram[15'h924] = 8'h06;
		ram[15'h925] = 8'h05;
		ram[15'h926] = 8'hCB;
		ram[15'h927] = 8'hE0;
		ram[15'h928] = 8'hCB;
		ram[15'h929] = 8'hE1;
		ram[15'h92A] = 8'hCB;
		ram[15'h92B] = 8'hE2;
		ram[15'h92C] = 8'hCB;
		ram[15'h92D] = 8'hE3;
		ram[15'h92E] = 8'hCB;
		ram[15'h92F] = 8'hE4;
		ram[15'h930] = 8'hCB;
		ram[15'h931] = 8'hE5;
		ram[15'h932] = 8'hCB;
		ram[15'h933] = 8'hE7;
		ram[15'h934] = 8'h21;
		ram[15'h935] = 8'h96;
		ram[15'h936] = 8'h00;
		ram[15'h937] = 8'hCB;
		ram[15'h938] = 8'hE6;
		ram[15'h939] = 8'hDD;
		ram[15'h93A] = 8'hCB;
		ram[15'h93B] = 8'h01;
		ram[15'h93C] = 8'hE6;
		ram[15'h93D] = 8'hFD;
		ram[15'h93E] = 8'hCB;
		ram[15'h93F] = 8'h02;
		ram[15'h940] = 8'hE6;
		ram[15'h941] = 8'h21;
		ram[15'h942] = 8'h06;
		ram[15'h943] = 8'h05;
		ram[15'h944] = 8'hCB;
		ram[15'h945] = 8'hA0;
		ram[15'h946] = 8'hCB;
		ram[15'h947] = 8'hA1;
		ram[15'h948] = 8'hCB;
		ram[15'h949] = 8'hA2;
		ram[15'h94A] = 8'hCB;
		ram[15'h94B] = 8'hA3;
		ram[15'h94C] = 8'hCB;
		ram[15'h94D] = 8'hA4;
		ram[15'h94E] = 8'hCB;
		ram[15'h94F] = 8'hA5;
		ram[15'h950] = 8'hCB;
		ram[15'h951] = 8'hA7;
		ram[15'h952] = 8'h21;
		ram[15'h953] = 8'h96;
		ram[15'h954] = 8'h00;
		ram[15'h955] = 8'hCB;
		ram[15'h956] = 8'hA6;
		ram[15'h957] = 8'hDD;
		ram[15'h958] = 8'hCB;
		ram[15'h959] = 8'h01;
		ram[15'h95A] = 8'hA6;
		ram[15'h95B] = 8'hFD;
		ram[15'h95C] = 8'hCB;
		ram[15'h95D] = 8'h02;
		ram[15'h95E] = 8'hA6;
		ram[15'h95F] = 8'h21;
		ram[15'h960] = 8'h06;
		ram[15'h961] = 8'h05;
		ram[15'h962] = 8'hCB;
		ram[15'h963] = 8'h68;
		ram[15'h964] = 8'hCB;
		ram[15'h965] = 8'h69;
		ram[15'h966] = 8'hCB;
		ram[15'h967] = 8'h6A;
		ram[15'h968] = 8'hCB;
		ram[15'h969] = 8'h6B;
		ram[15'h96A] = 8'hCB;
		ram[15'h96B] = 8'h6C;
		ram[15'h96C] = 8'hCB;
		ram[15'h96D] = 8'h6D;
		ram[15'h96E] = 8'hCB;
		ram[15'h96F] = 8'h6F;
		ram[15'h970] = 8'h21;
		ram[15'h971] = 8'h96;
		ram[15'h972] = 8'h00;
		ram[15'h973] = 8'hCB;
		ram[15'h974] = 8'h6E;
		ram[15'h975] = 8'hDD;
		ram[15'h976] = 8'hCB;
		ram[15'h977] = 8'h01;
		ram[15'h978] = 8'h6E;
		ram[15'h979] = 8'hFD;
		ram[15'h97A] = 8'hCB;
		ram[15'h97B] = 8'h02;
		ram[15'h97C] = 8'h6E;
		ram[15'h97D] = 8'h21;
		ram[15'h97E] = 8'h06;
		ram[15'h97F] = 8'h05;
		ram[15'h980] = 8'hCB;
		ram[15'h981] = 8'hE8;
		ram[15'h982] = 8'hCB;
		ram[15'h983] = 8'hE9;
		ram[15'h984] = 8'hCB;
		ram[15'h985] = 8'hEA;
		ram[15'h986] = 8'hCB;
		ram[15'h987] = 8'hEB;
		ram[15'h988] = 8'hCB;
		ram[15'h989] = 8'hEC;
		ram[15'h98A] = 8'hCB;
		ram[15'h98B] = 8'hED;
		ram[15'h98C] = 8'hCB;
		ram[15'h98D] = 8'hEF;
		ram[15'h98E] = 8'h21;
		ram[15'h98F] = 8'h96;
		ram[15'h990] = 8'h00;
		ram[15'h991] = 8'hCB;
		ram[15'h992] = 8'hEE;
		ram[15'h993] = 8'hDD;
		ram[15'h994] = 8'hCB;
		ram[15'h995] = 8'h01;
		ram[15'h996] = 8'hEE;
		ram[15'h997] = 8'hFD;
		ram[15'h998] = 8'hCB;
		ram[15'h999] = 8'h02;
		ram[15'h99A] = 8'hEE;
		ram[15'h99B] = 8'h21;
		ram[15'h99C] = 8'h06;
		ram[15'h99D] = 8'h05;
		ram[15'h99E] = 8'hCB;
		ram[15'h99F] = 8'hA8;
		ram[15'h9A0] = 8'hCB;
		ram[15'h9A1] = 8'hA9;
		ram[15'h9A2] = 8'hCB;
		ram[15'h9A3] = 8'hAA;
		ram[15'h9A4] = 8'hCB;
		ram[15'h9A5] = 8'hAB;
		ram[15'h9A6] = 8'hCB;
		ram[15'h9A7] = 8'hAC;
		ram[15'h9A8] = 8'hCB;
		ram[15'h9A9] = 8'hAD;
		ram[15'h9AA] = 8'hCB;
		ram[15'h9AB] = 8'hAF;
		ram[15'h9AC] = 8'h21;
		ram[15'h9AD] = 8'h96;
		ram[15'h9AE] = 8'h00;
		ram[15'h9AF] = 8'hCB;
		ram[15'h9B0] = 8'hAE;
		ram[15'h9B1] = 8'hDD;
		ram[15'h9B2] = 8'hCB;
		ram[15'h9B3] = 8'h01;
		ram[15'h9B4] = 8'hAE;
		ram[15'h9B5] = 8'hFD;
		ram[15'h9B6] = 8'hCB;
		ram[15'h9B7] = 8'h02;
		ram[15'h9B8] = 8'hAE;
		ram[15'h9B9] = 8'h21;
		ram[15'h9BA] = 8'h06;
		ram[15'h9BB] = 8'h05;
		ram[15'h9BC] = 8'hCB;
		ram[15'h9BD] = 8'h70;
		ram[15'h9BE] = 8'hCB;
		ram[15'h9BF] = 8'h71;
		ram[15'h9C0] = 8'hCB;
		ram[15'h9C1] = 8'h72;
		ram[15'h9C2] = 8'hCB;
		ram[15'h9C3] = 8'h73;
		ram[15'h9C4] = 8'hCB;
		ram[15'h9C5] = 8'h74;
		ram[15'h9C6] = 8'hCB;
		ram[15'h9C7] = 8'h75;
		ram[15'h9C8] = 8'hCB;
		ram[15'h9C9] = 8'h77;
		ram[15'h9CA] = 8'h21;
		ram[15'h9CB] = 8'h96;
		ram[15'h9CC] = 8'h00;
		ram[15'h9CD] = 8'hCB;
		ram[15'h9CE] = 8'h76;
		ram[15'h9CF] = 8'hDD;
		ram[15'h9D0] = 8'hCB;
		ram[15'h9D1] = 8'h01;
		ram[15'h9D2] = 8'h76;
		ram[15'h9D3] = 8'hFD;
		ram[15'h9D4] = 8'hCB;
		ram[15'h9D5] = 8'h02;
		ram[15'h9D6] = 8'h76;
		ram[15'h9D7] = 8'h21;
		ram[15'h9D8] = 8'h06;
		ram[15'h9D9] = 8'h05;
		ram[15'h9DA] = 8'hCB;
		ram[15'h9DB] = 8'hF0;
		ram[15'h9DC] = 8'hCB;
		ram[15'h9DD] = 8'hF1;
		ram[15'h9DE] = 8'hCB;
		ram[15'h9DF] = 8'hF2;
		ram[15'h9E0] = 8'hCB;
		ram[15'h9E1] = 8'hF3;
		ram[15'h9E2] = 8'hCB;
		ram[15'h9E3] = 8'hF4;
		ram[15'h9E4] = 8'hCB;
		ram[15'h9E5] = 8'hF5;
		ram[15'h9E6] = 8'hCB;
		ram[15'h9E7] = 8'hF7;
		ram[15'h9E8] = 8'h21;
		ram[15'h9E9] = 8'h96;
		ram[15'h9EA] = 8'h00;
		ram[15'h9EB] = 8'hCB;
		ram[15'h9EC] = 8'hF6;
		ram[15'h9ED] = 8'hDD;
		ram[15'h9EE] = 8'hCB;
		ram[15'h9EF] = 8'h01;
		ram[15'h9F0] = 8'hF6;
		ram[15'h9F1] = 8'hFD;
		ram[15'h9F2] = 8'hCB;
		ram[15'h9F3] = 8'h02;
		ram[15'h9F4] = 8'hF6;
		ram[15'h9F5] = 8'h21;
		ram[15'h9F6] = 8'h06;
		ram[15'h9F7] = 8'h05;
		ram[15'h9F8] = 8'hCB;
		ram[15'h9F9] = 8'hB0;
		ram[15'h9FA] = 8'hCB;
		ram[15'h9FB] = 8'hB1;
		ram[15'h9FC] = 8'hCB;
		ram[15'h9FD] = 8'hB2;
		ram[15'h9FE] = 8'hCB;
		ram[15'h9FF] = 8'hB3;
		ram[15'hA00] = 8'hCB;
		ram[15'hA01] = 8'hB4;
		ram[15'hA02] = 8'hCB;
		ram[15'hA03] = 8'hB5;
		ram[15'hA04] = 8'hCB;
		ram[15'hA05] = 8'hB7;
		ram[15'hA06] = 8'h21;
		ram[15'hA07] = 8'h96;
		ram[15'hA08] = 8'h00;
		ram[15'hA09] = 8'hCB;
		ram[15'hA0A] = 8'hB6;
		ram[15'hA0B] = 8'hDD;
		ram[15'hA0C] = 8'hCB;
		ram[15'hA0D] = 8'h01;
		ram[15'hA0E] = 8'hB6;
		ram[15'hA0F] = 8'hFD;
		ram[15'hA10] = 8'hCB;
		ram[15'hA11] = 8'h02;
		ram[15'hA12] = 8'hB6;
		ram[15'hA13] = 8'h21;
		ram[15'hA14] = 8'h06;
		ram[15'hA15] = 8'h05;
		ram[15'hA16] = 8'hCB;
		ram[15'hA17] = 8'h78;
		ram[15'hA18] = 8'hCB;
		ram[15'hA19] = 8'h79;
		ram[15'hA1A] = 8'hCB;
		ram[15'hA1B] = 8'h7A;
		ram[15'hA1C] = 8'hCB;
		ram[15'hA1D] = 8'h7B;
		ram[15'hA1E] = 8'hCB;
		ram[15'hA1F] = 8'h7C;
		ram[15'hA20] = 8'hCB;
		ram[15'hA21] = 8'h7D;
		ram[15'hA22] = 8'hCB;
		ram[15'hA23] = 8'h7F;
		ram[15'hA24] = 8'h21;
		ram[15'hA25] = 8'h96;
		ram[15'hA26] = 8'h00;
		ram[15'hA27] = 8'hCB;
		ram[15'hA28] = 8'h7E;
		ram[15'hA29] = 8'hDD;
		ram[15'hA2A] = 8'hCB;
		ram[15'hA2B] = 8'h01;
		ram[15'hA2C] = 8'h7E;
		ram[15'hA2D] = 8'hFD;
		ram[15'hA2E] = 8'hCB;
		ram[15'hA2F] = 8'h02;
		ram[15'hA30] = 8'h7E;
		ram[15'hA31] = 8'h21;
		ram[15'hA32] = 8'h06;
		ram[15'hA33] = 8'h05;
		ram[15'hA34] = 8'hCB;
		ram[15'hA35] = 8'hF8;
		ram[15'hA36] = 8'hCB;
		ram[15'hA37] = 8'hF9;
		ram[15'hA38] = 8'hCB;
		ram[15'hA39] = 8'hFA;
		ram[15'hA3A] = 8'hCB;
		ram[15'hA3B] = 8'hFB;
		ram[15'hA3C] = 8'hCB;
		ram[15'hA3D] = 8'hFC;
		ram[15'hA3E] = 8'hCB;
		ram[15'hA3F] = 8'hFD;
		ram[15'hA40] = 8'hCB;
		ram[15'hA41] = 8'hFF;
		ram[15'hA42] = 8'h21;
		ram[15'hA43] = 8'h96;
		ram[15'hA44] = 8'h00;
		ram[15'hA45] = 8'hCB;
		ram[15'hA46] = 8'hFE;
		ram[15'hA47] = 8'hDD;
		ram[15'hA48] = 8'hCB;
		ram[15'hA49] = 8'h01;
		ram[15'hA4A] = 8'hFE;
		ram[15'hA4B] = 8'hFD;
		ram[15'hA4C] = 8'hCB;
		ram[15'hA4D] = 8'h02;
		ram[15'hA4E] = 8'hFE;
		ram[15'hA4F] = 8'h21;
		ram[15'hA50] = 8'h06;
		ram[15'hA51] = 8'h05;
		ram[15'hA52] = 8'hCB;
		ram[15'hA53] = 8'hB8;
		ram[15'hA54] = 8'hCB;
		ram[15'hA55] = 8'hB9;
		ram[15'hA56] = 8'hCB;
		ram[15'hA57] = 8'hBA;
		ram[15'hA58] = 8'hCB;
		ram[15'hA59] = 8'hBB;
		ram[15'hA5A] = 8'hCB;
		ram[15'hA5B] = 8'hBC;
		ram[15'hA5C] = 8'hCB;
		ram[15'hA5D] = 8'hBD;
		ram[15'hA5E] = 8'hCB;
		ram[15'hA5F] = 8'hBF;
		ram[15'hA60] = 8'h21;
		ram[15'hA61] = 8'h96;
		ram[15'hA62] = 8'h00;
		ram[15'hA63] = 8'hCB;
		ram[15'hA64] = 8'hBE;
		ram[15'hA65] = 8'hDD;
		ram[15'hA66] = 8'hCB;
		ram[15'hA67] = 8'h01;
		ram[15'hA68] = 8'hBE;
		ram[15'hA69] = 8'hFD;
		ram[15'hA6A] = 8'hCB;
		ram[15'hA6B] = 8'h02;
		ram[15'hA6C] = 8'hBE;
		ram[15'hA6D] = 8'hC9;
		ram[15'hA6E] = 8'h3E;
		ram[15'hA6F] = 8'h0F;
		ram[15'hA70] = 8'hD3;
		ram[15'hA71] = 8'h01;
		ram[15'hA72] = 8'hC3;
		ram[15'hA73] = 8'h76;
		ram[15'hA74] = 8'h0A;
		ram[15'hA75] = 8'h00;
		ram[15'hA76] = 8'h18;
		ram[15'hA77] = 8'h01;
		ram[15'hA78] = 8'h00;
		ram[15'hA79] = 8'hF3;
		ram[15'hA7A] = 8'h21;
		ram[15'hA7B] = 8'h00;
		ram[15'hA7C] = 8'h00;
		ram[15'hA7D] = 8'hE5;
		ram[15'hA7E] = 8'hF1;
		ram[15'hA7F] = 8'hCA;
		ram[15'hA80] = 8'hDB;
		ram[15'hA81] = 8'h0B;
		ram[15'hA82] = 8'hC2;
		ram[15'hA83] = 8'h86;
		ram[15'hA84] = 8'h0A;
		ram[15'hA85] = 8'h76;
		ram[15'hA86] = 8'hDA;
		ram[15'hA87] = 8'hDB;
		ram[15'hA88] = 8'h0B;
		ram[15'hA89] = 8'hD2;
		ram[15'hA8A] = 8'h8D;
		ram[15'hA8B] = 8'h0A;
		ram[15'hA8C] = 8'h76;
		ram[15'hA8D] = 8'hEA;
		ram[15'hA8E] = 8'hDB;
		ram[15'hA8F] = 8'h0B;
		ram[15'hA90] = 8'hE2;
		ram[15'hA91] = 8'h94;
		ram[15'hA92] = 8'h0A;
		ram[15'hA93] = 8'h76;
		ram[15'hA94] = 8'hFA;
		ram[15'hA95] = 8'hDB;
		ram[15'hA96] = 8'h0B;
		ram[15'hA97] = 8'hF2;
		ram[15'hA98] = 8'h9B;
		ram[15'hA99] = 8'h0A;
		ram[15'hA9A] = 8'h76;
		ram[15'hA9B] = 8'h21;
		ram[15'hA9C] = 8'h01;
		ram[15'hA9D] = 8'h00;
		ram[15'hA9E] = 8'hE5;
		ram[15'hA9F] = 8'hF1;
		ram[15'hAA0] = 8'hD2;
		ram[15'hAA1] = 8'hDB;
		ram[15'hAA2] = 8'h0B;
		ram[15'hAA3] = 8'hDA;
		ram[15'hAA4] = 8'hA7;
		ram[15'hAA5] = 8'h0A;
		ram[15'hAA6] = 8'h76;
		ram[15'hAA7] = 8'h21;
		ram[15'hAA8] = 8'h40;
		ram[15'hAA9] = 8'h00;
		ram[15'hAAA] = 8'hE5;
		ram[15'hAAB] = 8'hF1;
		ram[15'hAAC] = 8'hC2;
		ram[15'hAAD] = 8'hDB;
		ram[15'hAAE] = 8'h0B;
		ram[15'hAAF] = 8'hCA;
		ram[15'hAB0] = 8'hB3;
		ram[15'hAB1] = 8'h0A;
		ram[15'hAB2] = 8'h76;
		ram[15'hAB3] = 8'h21;
		ram[15'hAB4] = 8'h04;
		ram[15'hAB5] = 8'h00;
		ram[15'hAB6] = 8'hE5;
		ram[15'hAB7] = 8'hF1;
		ram[15'hAB8] = 8'hE2;
		ram[15'hAB9] = 8'hDB;
		ram[15'hABA] = 8'h0B;
		ram[15'hABB] = 8'hEA;
		ram[15'hABC] = 8'hBF;
		ram[15'hABD] = 8'h0A;
		ram[15'hABE] = 8'h76;
		ram[15'hABF] = 8'h21;
		ram[15'hAC0] = 8'h80;
		ram[15'hAC1] = 8'h00;
		ram[15'hAC2] = 8'hE5;
		ram[15'hAC3] = 8'hF1;
		ram[15'hAC4] = 8'hF2;
		ram[15'hAC5] = 8'hDB;
		ram[15'hAC6] = 8'h0B;
		ram[15'hAC7] = 8'hFA;
		ram[15'hAC8] = 8'hCB;
		ram[15'hAC9] = 8'h0A;
		ram[15'hACA] = 8'h76;
		ram[15'hACB] = 8'h21;
		ram[15'hACC] = 8'h00;
		ram[15'hACD] = 8'h00;
		ram[15'hACE] = 8'hE5;
		ram[15'hACF] = 8'hF1;
		ram[15'hAD0] = 8'h38;
		ram[15'hAD1] = 8'h02;
		ram[15'hAD2] = 8'h30;
		ram[15'hAD3] = 8'h01;
		ram[15'hAD4] = 8'h76;
		ram[15'hAD5] = 8'h28;
		ram[15'hAD6] = 8'hFD;
		ram[15'hAD7] = 8'h20;
		ram[15'hAD8] = 8'h01;
		ram[15'hAD9] = 8'h76;
		ram[15'hADA] = 8'h21;
		ram[15'hADB] = 8'h40;
		ram[15'hADC] = 8'h00;
		ram[15'hADD] = 8'hE5;
		ram[15'hADE] = 8'hF1;
		ram[15'hADF] = 8'h20;
		ram[15'hAE0] = 8'hF3;
		ram[15'hAE1] = 8'h28;
		ram[15'hAE2] = 8'h01;
		ram[15'hAE3] = 8'h76;
		ram[15'hAE4] = 8'h21;
		ram[15'hAE5] = 8'h01;
		ram[15'hAE6] = 8'h00;
		ram[15'hAE7] = 8'hE5;
		ram[15'hAE8] = 8'hF1;
		ram[15'hAE9] = 8'h30;
		ram[15'hAEA] = 8'hE9;
		ram[15'hAEB] = 8'h38;
		ram[15'hAEC] = 8'h01;
		ram[15'hAED] = 8'h76;
		ram[15'hAEE] = 8'h21;
		ram[15'hAEF] = 8'hF2;
		ram[15'hAF0] = 8'h0A;
		ram[15'hAF1] = 8'hE9;
		ram[15'hAF2] = 8'hDD;
		ram[15'hAF3] = 8'h21;
		ram[15'hAF4] = 8'hF8;
		ram[15'hAF5] = 8'h0A;
		ram[15'hAF6] = 8'hDD;
		ram[15'hAF7] = 8'hE9;
		ram[15'hAF8] = 8'hFD;
		ram[15'hAF9] = 8'h21;
		ram[15'hAFA] = 8'hFE;
		ram[15'hAFB] = 8'h0A;
		ram[15'hAFC] = 8'hFD;
		ram[15'hAFD] = 8'hE9;
		ram[15'hAFE] = 8'h21;
		ram[15'hAFF] = 8'h92;
		ram[15'hB00] = 8'h00;
		ram[15'hB01] = 8'h01;
		ram[15'hB02] = 8'h00;
		ram[15'hB03] = 8'h05;
		ram[15'hB04] = 8'h70;
		ram[15'hB05] = 8'h10;
		ram[15'hB06] = 8'hFD;
		ram[15'hB07] = 8'hFB;
		ram[15'hB08] = 8'hC9;
		ram[15'hB09] = 8'hF3;
		ram[15'hB0A] = 8'h3E;
		ram[15'hB0B] = 8'h10;
		ram[15'hB0C] = 8'hD3;
		ram[15'hB0D] = 8'h01;
		ram[15'hB0E] = 8'h21;
		ram[15'hB0F] = 8'h00;
		ram[15'hB10] = 8'h00;
		ram[15'hB11] = 8'hE5;
		ram[15'hB12] = 8'hF1;
		ram[15'hB13] = 8'hDC;
		ram[15'hB14] = 8'hDB;
		ram[15'hB15] = 8'h0B;
		ram[15'hB16] = 8'hD4;
		ram[15'hB17] = 8'h1A;
		ram[15'hB18] = 8'h0B;
		ram[15'hB19] = 8'h76;
		ram[15'hB1A] = 8'hD1;
		ram[15'hB1B] = 8'hCC;
		ram[15'hB1C] = 8'hDB;
		ram[15'hB1D] = 8'h0B;
		ram[15'hB1E] = 8'hC4;
		ram[15'hB1F] = 8'h22;
		ram[15'hB20] = 8'h0B;
		ram[15'hB21] = 8'h76;
		ram[15'hB22] = 8'hD1;
		ram[15'hB23] = 8'hEC;
		ram[15'hB24] = 8'hDB;
		ram[15'hB25] = 8'h0B;
		ram[15'hB26] = 8'hE4;
		ram[15'hB27] = 8'h2A;
		ram[15'hB28] = 8'h0B;
		ram[15'hB29] = 8'h76;
		ram[15'hB2A] = 8'hD1;
		ram[15'hB2B] = 8'hFC;
		ram[15'hB2C] = 8'hDB;
		ram[15'hB2D] = 8'h0B;
		ram[15'hB2E] = 8'hF4;
		ram[15'hB2F] = 8'h32;
		ram[15'hB30] = 8'h0B;
		ram[15'hB31] = 8'h76;
		ram[15'hB32] = 8'hD1;
		ram[15'hB33] = 8'h21;
		ram[15'hB34] = 8'h01;
		ram[15'hB35] = 8'h00;
		ram[15'hB36] = 8'hE5;
		ram[15'hB37] = 8'hF1;
		ram[15'hB38] = 8'hD4;
		ram[15'hB39] = 8'hDB;
		ram[15'hB3A] = 8'h0B;
		ram[15'hB3B] = 8'hDC;
		ram[15'hB3C] = 8'h3F;
		ram[15'hB3D] = 8'h0B;
		ram[15'hB3E] = 8'h76;
		ram[15'hB3F] = 8'hD1;
		ram[15'hB40] = 8'h21;
		ram[15'hB41] = 8'h40;
		ram[15'hB42] = 8'h00;
		ram[15'hB43] = 8'hE5;
		ram[15'hB44] = 8'hF1;
		ram[15'hB45] = 8'hC4;
		ram[15'hB46] = 8'hDB;
		ram[15'hB47] = 8'h0B;
		ram[15'hB48] = 8'hCC;
		ram[15'hB49] = 8'h4C;
		ram[15'hB4A] = 8'h0B;
		ram[15'hB4B] = 8'h76;
		ram[15'hB4C] = 8'hD1;
		ram[15'hB4D] = 8'h21;
		ram[15'hB4E] = 8'h04;
		ram[15'hB4F] = 8'h00;
		ram[15'hB50] = 8'hE5;
		ram[15'hB51] = 8'hF1;
		ram[15'hB52] = 8'hE4;
		ram[15'hB53] = 8'hDB;
		ram[15'hB54] = 8'h0B;
		ram[15'hB55] = 8'hEC;
		ram[15'hB56] = 8'h59;
		ram[15'hB57] = 8'h0B;
		ram[15'hB58] = 8'h76;
		ram[15'hB59] = 8'hD1;
		ram[15'hB5A] = 8'h21;
		ram[15'hB5B] = 8'h80;
		ram[15'hB5C] = 8'h00;
		ram[15'hB5D] = 8'hE5;
		ram[15'hB5E] = 8'hF1;
		ram[15'hB5F] = 8'hF4;
		ram[15'hB60] = 8'hDB;
		ram[15'hB61] = 8'h0B;
		ram[15'hB62] = 8'hFC;
		ram[15'hB63] = 8'h66;
		ram[15'hB64] = 8'h0B;
		ram[15'hB65] = 8'h76;
		ram[15'hB66] = 8'hD1;
		ram[15'hB67] = 8'h01;
		ram[15'hB68] = 8'hDB;
		ram[15'hB69] = 8'h0B;
		ram[15'hB6A] = 8'h21;
		ram[15'hB6B] = 8'h00;
		ram[15'hB6C] = 8'h00;
		ram[15'hB6D] = 8'hE5;
		ram[15'hB6E] = 8'hF1;
		ram[15'hB6F] = 8'hC5;
		ram[15'hB70] = 8'hD8;
		ram[15'hB71] = 8'hC1;
		ram[15'hB72] = 8'h21;
		ram[15'hB73] = 8'h78;
		ram[15'hB74] = 8'h0B;
		ram[15'hB75] = 8'hE5;
		ram[15'hB76] = 8'hD0;
		ram[15'hB77] = 8'h76;
		ram[15'hB78] = 8'hC5;
		ram[15'hB79] = 8'hC8;
		ram[15'hB7A] = 8'hC1;
		ram[15'hB7B] = 8'h21;
		ram[15'hB7C] = 8'h81;
		ram[15'hB7D] = 8'h0B;
		ram[15'hB7E] = 8'hE5;
		ram[15'hB7F] = 8'hC0;
		ram[15'hB80] = 8'h76;
		ram[15'hB81] = 8'hC5;
		ram[15'hB82] = 8'hE8;
		ram[15'hB83] = 8'hC1;
		ram[15'hB84] = 8'h21;
		ram[15'hB85] = 8'h8A;
		ram[15'hB86] = 8'h0B;
		ram[15'hB87] = 8'hE5;
		ram[15'hB88] = 8'hE0;
		ram[15'hB89] = 8'h76;
		ram[15'hB8A] = 8'hC5;
		ram[15'hB8B] = 8'hF8;
		ram[15'hB8C] = 8'hC1;
		ram[15'hB8D] = 8'h21;
		ram[15'hB8E] = 8'h93;
		ram[15'hB8F] = 8'h0B;
		ram[15'hB90] = 8'hE5;
		ram[15'hB91] = 8'hF0;
		ram[15'hB92] = 8'h76;
		ram[15'hB93] = 8'h21;
		ram[15'hB94] = 8'h01;
		ram[15'hB95] = 8'h00;
		ram[15'hB96] = 8'hE5;
		ram[15'hB97] = 8'hF1;
		ram[15'hB98] = 8'hC5;
		ram[15'hB99] = 8'hD0;
		ram[15'hB9A] = 8'hC1;
		ram[15'hB9B] = 8'h21;
		ram[15'hB9C] = 8'hA1;
		ram[15'hB9D] = 8'h0B;
		ram[15'hB9E] = 8'hE5;
		ram[15'hB9F] = 8'hD8;
		ram[15'hBA0] = 8'h76;
		ram[15'hBA1] = 8'h21;
		ram[15'hBA2] = 8'h40;
		ram[15'hBA3] = 8'h00;
		ram[15'hBA4] = 8'hE5;
		ram[15'hBA5] = 8'hF1;
		ram[15'hBA6] = 8'hC5;
		ram[15'hBA7] = 8'hC0;
		ram[15'hBA8] = 8'hC1;
		ram[15'hBA9] = 8'h21;
		ram[15'hBAA] = 8'hAF;
		ram[15'hBAB] = 8'h0B;
		ram[15'hBAC] = 8'hE5;
		ram[15'hBAD] = 8'hC8;
		ram[15'hBAE] = 8'h76;
		ram[15'hBAF] = 8'h21;
		ram[15'hBB0] = 8'h04;
		ram[15'hBB1] = 8'h00;
		ram[15'hBB2] = 8'hE5;
		ram[15'hBB3] = 8'hF1;
		ram[15'hBB4] = 8'hC5;
		ram[15'hBB5] = 8'hE0;
		ram[15'hBB6] = 8'hC1;
		ram[15'hBB7] = 8'h21;
		ram[15'hBB8] = 8'hBD;
		ram[15'hBB9] = 8'h0B;
		ram[15'hBBA] = 8'hE5;
		ram[15'hBBB] = 8'hE8;
		ram[15'hBBC] = 8'h76;
		ram[15'hBBD] = 8'h21;
		ram[15'hBBE] = 8'h80;
		ram[15'hBBF] = 8'h00;
		ram[15'hBC0] = 8'hE5;
		ram[15'hBC1] = 8'hF1;
		ram[15'hBC2] = 8'hC5;
		ram[15'hBC3] = 8'hF0;
		ram[15'hBC4] = 8'hC1;
		ram[15'hBC5] = 8'h21;
		ram[15'hBC6] = 8'hCB;
		ram[15'hBC7] = 8'h0B;
		ram[15'hBC8] = 8'hE5;
		ram[15'hBC9] = 8'hF8;
		ram[15'hBCA] = 8'h76;
		ram[15'hBCB] = 8'hCD;
		ram[15'hBCC] = 8'hCF;
		ram[15'hBCD] = 8'h0B;
		ram[15'hBCE] = 8'h76;
		ram[15'hBCF] = 8'hD1;
		ram[15'hBD0] = 8'h21;
		ram[15'hBD1] = 8'hD9;
		ram[15'hBD2] = 8'h0B;
		ram[15'hBD3] = 8'hE5;
		ram[15'hBD4] = 8'hC9;
		ram[15'hBD5] = 8'h76;
		ram[15'hBD6] = 8'hDF;
		ram[15'hBD7] = 8'hE7;
		ram[15'hBD8] = 8'hEF;
		ram[15'hBD9] = 8'hFB;
		ram[15'hBDA] = 8'hC9;
		ram[15'hBDB] = 8'h76;
		ram[15'hBDC] = 8'h3E;
		ram[15'hBDD] = 8'h11;
		ram[15'hBDE] = 8'hD3;
		ram[15'hBDF] = 8'h01;
		ram[15'hBE0] = 8'h3E;
		ram[15'hBE1] = 8'h00;
		ram[15'hBE2] = 8'hDB;
		ram[15'hBE3] = 8'h02;
		ram[15'hBE4] = 8'h32;
		ram[15'hBE5] = 8'h92;
		ram[15'hBE6] = 8'h00;
		ram[15'hBE7] = 8'h01;
		ram[15'hBE8] = 8'h03;
		ram[15'hBE9] = 8'h00;
		ram[15'hBEA] = 8'hED;
		ram[15'hBEB] = 8'h78;
		ram[15'hBEC] = 8'hED;
		ram[15'hBED] = 8'h50;
		ram[15'hBEE] = 8'hED;
		ram[15'hBEF] = 8'h58;
		ram[15'hBF0] = 8'hED;
		ram[15'hBF1] = 8'h60;
		ram[15'hBF2] = 8'hED;
		ram[15'hBF3] = 8'h68;
		ram[15'hBF4] = 8'hED;
		ram[15'hBF5] = 8'h40;
		ram[15'hBF6] = 8'h06;
		ram[15'hBF7] = 8'h00;
		ram[15'hBF8] = 8'hED;
		ram[15'hBF9] = 8'h48;
		ram[15'hBFA] = 8'h3E;
		ram[15'hBFB] = 8'h55;
		ram[15'hBFC] = 8'hD3;
		ram[15'hBFD] = 8'h02;
		ram[15'hBFE] = 8'h01;
		ram[15'hBFF] = 8'h03;
		ram[15'hC00] = 8'h00;
		ram[15'hC01] = 8'h11;
		ram[15'hC02] = 8'h05;
		ram[15'hC03] = 8'h04;
		ram[15'hC04] = 8'h21;
		ram[15'hC05] = 8'h07;
		ram[15'hC06] = 8'h06;
		ram[15'hC07] = 8'hED;
		ram[15'hC08] = 8'h41;
		ram[15'hC09] = 8'hED;
		ram[15'hC0A] = 8'h49;
		ram[15'hC0B] = 8'hED;
		ram[15'hC0C] = 8'h51;
		ram[15'hC0D] = 8'hED;
		ram[15'hC0E] = 8'h59;
		ram[15'hC0F] = 8'hED;
		ram[15'hC10] = 8'h61;
		ram[15'hC11] = 8'hED;
		ram[15'hC12] = 8'h69;
		ram[15'hC13] = 8'h21;
		ram[15'hC14] = 8'h98;
		ram[15'hC15] = 8'h00;
		ram[15'hC16] = 8'h01;
		ram[15'hC17] = 8'hFF;
		ram[15'hC18] = 8'h01;
		ram[15'hC19] = 8'hED;
		ram[15'hC1A] = 8'hA2;
		ram[15'hC1B] = 8'hED;
		ram[15'hC1C] = 8'hA2;
		ram[15'hC1D] = 8'hED;
		ram[15'hC1E] = 8'hA2;
		ram[15'hC1F] = 8'hED;
		ram[15'hC20] = 8'hA2;
		ram[15'hC21] = 8'h22;
		ram[15'hC22] = 8'h96;
		ram[15'hC23] = 8'h00;
		ram[15'hC24] = 8'hED;
		ram[15'hC25] = 8'h43;
		ram[15'hC26] = 8'h96;
		ram[15'hC27] = 8'h00;
		ram[15'hC28] = 8'h21;
		ram[15'hC29] = 8'hA7;
		ram[15'hC2A] = 8'h00;
		ram[15'hC2B] = 8'h01;
		ram[15'hC2C] = 8'hFF;
		ram[15'hC2D] = 8'h01;
		ram[15'hC2E] = 8'hED;
		ram[15'hC2F] = 8'hAA;
		ram[15'hC30] = 8'hED;
		ram[15'hC31] = 8'hAA;
		ram[15'hC32] = 8'hED;
		ram[15'hC33] = 8'hAA;
		ram[15'hC34] = 8'hED;
		ram[15'hC35] = 8'hAA;
		ram[15'hC36] = 8'h22;
		ram[15'hC37] = 8'h96;
		ram[15'hC38] = 8'h00;
		ram[15'hC39] = 8'hED;
		ram[15'hC3A] = 8'h43;
		ram[15'hC3B] = 8'h96;
		ram[15'hC3C] = 8'h00;
		ram[15'hC3D] = 8'h21;
		ram[15'hC3E] = 8'h98;
		ram[15'hC3F] = 8'h00;
		ram[15'hC40] = 8'h01;
		ram[15'hC41] = 8'hFF;
		ram[15'hC42] = 8'h01;
		ram[15'hC43] = 8'hED;
		ram[15'hC44] = 8'hA3;
		ram[15'hC45] = 8'hED;
		ram[15'hC46] = 8'hA3;
		ram[15'hC47] = 8'hED;
		ram[15'hC48] = 8'hA3;
		ram[15'hC49] = 8'hED;
		ram[15'hC4A] = 8'hA3;
		ram[15'hC4B] = 8'h22;
		ram[15'hC4C] = 8'h96;
		ram[15'hC4D] = 8'h00;
		ram[15'hC4E] = 8'hED;
		ram[15'hC4F] = 8'h43;
		ram[15'hC50] = 8'h96;
		ram[15'hC51] = 8'h00;
		ram[15'hC52] = 8'h21;
		ram[15'hC53] = 8'hA7;
		ram[15'hC54] = 8'h00;
		ram[15'hC55] = 8'h01;
		ram[15'hC56] = 8'hFF;
		ram[15'hC57] = 8'h01;
		ram[15'hC58] = 8'hED;
		ram[15'hC59] = 8'hAB;
		ram[15'hC5A] = 8'hED;
		ram[15'hC5B] = 8'hAB;
		ram[15'hC5C] = 8'hED;
		ram[15'hC5D] = 8'hAB;
		ram[15'hC5E] = 8'hED;
		ram[15'hC5F] = 8'hAB;
		ram[15'hC60] = 8'h22;
		ram[15'hC61] = 8'h96;
		ram[15'hC62] = 8'h00;
		ram[15'hC63] = 8'hED;
		ram[15'hC64] = 8'h43;
		ram[15'hC65] = 8'h96;
		ram[15'hC66] = 8'h00;
		ram[15'hC67] = 8'h21;
		ram[15'hC68] = 8'h98;
		ram[15'hC69] = 8'h00;
		ram[15'hC6A] = 8'h01;
		ram[15'hC6B] = 8'hFF;
		ram[15'hC6C] = 8'h05;
		ram[15'hC6D] = 8'hED;
		ram[15'hC6E] = 8'hB2;
		ram[15'hC6F] = 8'h22;
		ram[15'hC70] = 8'h96;
		ram[15'hC71] = 8'h00;
		ram[15'hC72] = 8'hED;
		ram[15'hC73] = 8'h43;
		ram[15'hC74] = 8'h96;
		ram[15'hC75] = 8'h00;
		ram[15'hC76] = 8'h21;
		ram[15'hC77] = 8'hA7;
		ram[15'hC78] = 8'h00;
		ram[15'hC79] = 8'h01;
		ram[15'hC7A] = 8'hFF;
		ram[15'hC7B] = 8'h05;
		ram[15'hC7C] = 8'hED;
		ram[15'hC7D] = 8'hB2;
		ram[15'hC7E] = 8'h22;
		ram[15'hC7F] = 8'h96;
		ram[15'hC80] = 8'h00;
		ram[15'hC81] = 8'hED;
		ram[15'hC82] = 8'h43;
		ram[15'hC83] = 8'h96;
		ram[15'hC84] = 8'h00;
		ram[15'hC85] = 8'h21;
		ram[15'hC86] = 8'h98;
		ram[15'hC87] = 8'h00;
		ram[15'hC88] = 8'h01;
		ram[15'hC89] = 8'hFF;
		ram[15'hC8A] = 8'h05;
		ram[15'hC8B] = 8'hED;
		ram[15'hC8C] = 8'hB3;
		ram[15'hC8D] = 8'h22;
		ram[15'hC8E] = 8'h96;
		ram[15'hC8F] = 8'h00;
		ram[15'hC90] = 8'hED;
		ram[15'hC91] = 8'h43;
		ram[15'hC92] = 8'h96;
		ram[15'hC93] = 8'h00;
		ram[15'hC94] = 8'h21;
		ram[15'hC95] = 8'hA7;
		ram[15'hC96] = 8'h00;
		ram[15'hC97] = 8'h01;
		ram[15'hC98] = 8'hFF;
		ram[15'hC99] = 8'h05;
		ram[15'hC9A] = 8'hED;
		ram[15'hC9B] = 8'hBB;
		ram[15'hC9C] = 8'h22;
		ram[15'hC9D] = 8'h96;
		ram[15'hC9E] = 8'h00;
		ram[15'hC9F] = 8'hED;
		ram[15'hCA0] = 8'h43;
		ram[15'hCA1] = 8'h96;
		ram[15'hCA2] = 8'h00;
		ram[15'hCA3] = 8'hC9;
		ram[15'hCA4] = 8'hF5;
		ram[15'hCA5] = 8'hC5;
		ram[15'hCA6] = 8'hD5;
		ram[15'hCA7] = 8'hE5;
		ram[15'hCA8] = 8'h47;
		ram[15'hCA9] = 8'h79;
		ram[15'hCAA] = 8'hFE;
		ram[15'hCAB] = 8'h02;
		ram[15'hCAC] = 8'h28;
		ram[15'hCAD] = 8'h09;
		ram[15'hCAE] = 8'hFE;
		ram[15'hCAF] = 8'h09;
		ram[15'hCB0] = 8'h28;
		ram[15'hCB1] = 8'h0D;
		ram[15'hCB2] = 8'hE1;
		ram[15'hCB3] = 8'hD1;
		ram[15'hCB4] = 8'hC1;
		ram[15'hCB5] = 8'hF1;
		ram[15'hCB6] = 8'hC9;
		ram[15'hCB7] = 8'h78;
		ram[15'hCB8] = 8'hFE;
		ram[15'hCB9] = 8'h0A;
		ram[15'hCBA] = 8'h28;
		ram[15'hCBB] = 8'hF6;
		ram[15'hCBC] = 8'hD7;
		ram[15'hCBD] = 8'h18;
		ram[15'hCBE] = 8'hF3;
		ram[15'hCBF] = 8'h1A;
		ram[15'hCC0] = 8'hFE;
		ram[15'hCC1] = 8'h00;
		ram[15'hCC2] = 8'h28;
		ram[15'hCC3] = 8'hEE;
		ram[15'hCC4] = 8'hFE;
		ram[15'hCC5] = 8'h0A;
		ram[15'hCC6] = 8'hC4;
		ram[15'hCC7] = 8'h10;
		ram[15'hCC8] = 8'h00;
		ram[15'hCC9] = 8'h13;
		ram[15'hCCA] = 8'h18;
		ram[15'hCCB] = 8'hF3;
		ram[15'hCCC] = 8'h00;
		ram[15'hCCD] = 8'h00;
		ram[15'hCCE] = 8'h00;
		ram[15'hCCF] = 8'h00;
		ram[15'hCD0] = 8'h00;
		ram[15'hCD1] = 8'h00;
		ram[15'hCD2] = 8'h00;
		ram[15'hCD3] = 8'h00;
		ram[15'hCD4] = 8'h00;
		ram[15'hCD5] = 8'h00;
		ram[15'hCD6] = 8'h00;
		ram[15'hCD7] = 8'h00;
		ram[15'hCD8] = 8'h00;
		ram[15'hCD9] = 8'h00;
		ram[15'hCDA] = 8'h00;
		ram[15'hCDB] = 8'h00;
		ram[15'hCDC] = 8'h00;
		ram[15'hCDD] = 8'h00;
		ram[15'hCDE] = 8'h00;
		ram[15'hCDF] = 8'h00;
		ram[15'hCE0] = 8'h00;
		ram[15'hCE1] = 8'h00;
		ram[15'hCE2] = 8'h00;
		ram[15'hCE3] = 8'h00;
		ram[15'hCE4] = 8'h00;
		ram[15'hCE5] = 8'h00;
		ram[15'hCE6] = 8'h00;
		ram[15'hCE7] = 8'h00;
		ram[15'hCE8] = 8'h00;
		ram[15'hCE9] = 8'h00;
		ram[15'hCEA] = 8'h00;
		ram[15'hCEB] = 8'h00;


		
end

endmodule 